/*  This module contains the codepage 437 font ROM.
*/
module font437(clk, char, row, bits);
    input clk;           // clock
    input [7:0] char;    // character to display
    input [3:0] row;     // font row # in char
    output [7:0] bits;   // output (8 bits)

    // font array (256 x 12 x 8 bits)
    reg   [7:0] font437[3071:0];
    reg   [7:0] fontrow; // row of data from font
    wire  [11:0] faddr;  // address in font array

    initial begin
        font437[0] = 8'b00000000;
        font437[1] = 8'b00000000;
        font437[2] = 8'b00000000;
        font437[3] = 8'b00000000;
        font437[4] = 8'b00000000;
        font437[5] = 8'b00000000;
        font437[6] = 8'b00000000;
        font437[7] = 8'b00000000;
        font437[8] = 8'b00000000;
        font437[9] = 8'b00000000;
        font437[10] = 8'b00000000;
        font437[11] = 8'b00000000;
        font437[12] = 8'b00000000;
        font437[13] = 8'b01111110;
        font437[14] = 8'b11000011;
        font437[15] = 8'b10000001;
        font437[16] = 8'b10100101;
        font437[17] = 8'b10000001;
        font437[18] = 8'b10111101;
        font437[19] = 8'b10011001;
        font437[20] = 8'b11000011;
        font437[21] = 8'b01111110;
        font437[22] = 8'b00000000;
        font437[23] = 8'b00000000;
        font437[24] = 8'b00000000;
        font437[25] = 8'b01111110;
        font437[26] = 8'b11111111;
        font437[27] = 8'b11111111;
        font437[28] = 8'b11011011;
        font437[29] = 8'b11111111;
        font437[30] = 8'b11000011;
        font437[31] = 8'b11100111;
        font437[32] = 8'b11111111;
        font437[33] = 8'b01111110;
        font437[34] = 8'b00000000;
        font437[35] = 8'b00000000;
        font437[36] = 8'b00000000;
        font437[37] = 8'b00000000;
        font437[38] = 8'b01000100;
        font437[39] = 8'b11101110;
        font437[40] = 8'b11111110;
        font437[41] = 8'b11111110;
        font437[42] = 8'b11111110;
        font437[43] = 8'b01111100;
        font437[44] = 8'b00111000;
        font437[45] = 8'b00010000;
        font437[46] = 8'b00000000;
        font437[47] = 8'b00000000;
        font437[48] = 8'b00000000;
        font437[49] = 8'b00010000;
        font437[50] = 8'b00111000;
        font437[51] = 8'b01111100;
        font437[52] = 8'b11111110;
        font437[53] = 8'b11111110;
        font437[54] = 8'b01111100;
        font437[55] = 8'b00111000;
        font437[56] = 8'b00010000;
        font437[57] = 8'b00000000;
        font437[58] = 8'b00000000;
        font437[59] = 8'b00000000;
        font437[60] = 8'b00000000;
        font437[61] = 8'b00011000;
        font437[62] = 8'b00111100;
        font437[63] = 8'b00111100;
        font437[64] = 8'b11111111;
        font437[65] = 8'b11100111;
        font437[66] = 8'b11100111;
        font437[67] = 8'b00011000;
        font437[68] = 8'b00011000;
        font437[69] = 8'b01111110;
        font437[70] = 8'b00000000;
        font437[71] = 8'b00000000;
        font437[72] = 8'b00000000;
        font437[73] = 8'b00011000;
        font437[74] = 8'b00111100;
        font437[75] = 8'b01111110;
        font437[76] = 8'b11111111;
        font437[77] = 8'b11111111;
        font437[78] = 8'b01111110;
        font437[79] = 8'b00011000;
        font437[80] = 8'b00011000;
        font437[81] = 8'b01111110;
        font437[82] = 8'b00000000;
        font437[83] = 8'b00000000;
        font437[84] = 8'b00000000;
        font437[85] = 8'b00000000;
        font437[86] = 8'b00000000;
        font437[87] = 8'b00000000;
        font437[88] = 8'b00111100;
        font437[89] = 8'b01111110;
        font437[90] = 8'b01111110;
        font437[91] = 8'b00111100;
        font437[92] = 8'b00000000;
        font437[93] = 8'b00000000;
        font437[94] = 8'b00000000;
        font437[95] = 8'b00000000;
        font437[96] = 8'b11111111;
        font437[97] = 8'b11111111;
        font437[98] = 8'b11111111;
        font437[99] = 8'b11111111;
        font437[100] = 8'b11000011;
        font437[101] = 8'b10000001;
        font437[102] = 8'b10000001;
        font437[103] = 8'b11000011;
        font437[104] = 8'b11111111;
        font437[105] = 8'b11111111;
        font437[106] = 8'b11111111;
        font437[107] = 8'b11111111;
        font437[108] = 8'b00000000;
        font437[109] = 8'b00000000;
        font437[110] = 8'b00111100;
        font437[111] = 8'b01111110;
        font437[112] = 8'b01100110;
        font437[113] = 8'b01000010;
        font437[114] = 8'b01000010;
        font437[115] = 8'b01100110;
        font437[116] = 8'b01111110;
        font437[117] = 8'b00111100;
        font437[118] = 8'b00000000;
        font437[119] = 8'b00000000;
        font437[120] = 8'b11111111;
        font437[121] = 8'b11111111;
        font437[122] = 8'b11000011;
        font437[123] = 8'b10000001;
        font437[124] = 8'b10011001;
        font437[125] = 8'b10111101;
        font437[126] = 8'b10111101;
        font437[127] = 8'b10011001;
        font437[128] = 8'b10000001;
        font437[129] = 8'b11000011;
        font437[130] = 8'b11111111;
        font437[131] = 8'b11111111;
        font437[132] = 8'b00000000;
        font437[133] = 8'b00111110;
        font437[134] = 8'b00001110;
        font437[135] = 8'b00111010;
        font437[136] = 8'b01110010;
        font437[137] = 8'b11111000;
        font437[138] = 8'b11001100;
        font437[139] = 8'b11001100;
        font437[140] = 8'b11001100;
        font437[141] = 8'b01111000;
        font437[142] = 8'b00000000;
        font437[143] = 8'b00000000;
        font437[144] = 8'b00000000;
        font437[145] = 8'b00111100;
        font437[146] = 8'b01100110;
        font437[147] = 8'b01100110;
        font437[148] = 8'b01100110;
        font437[149] = 8'b00111100;
        font437[150] = 8'b00011000;
        font437[151] = 8'b01111110;
        font437[152] = 8'b00011000;
        font437[153] = 8'b00011000;
        font437[154] = 8'b00000000;
        font437[155] = 8'b00000000;
        font437[156] = 8'b00000000;
        font437[157] = 8'b00011111;
        font437[158] = 8'b00011001;
        font437[159] = 8'b00011001;
        font437[160] = 8'b00011111;
        font437[161] = 8'b00011000;
        font437[162] = 8'b00011000;
        font437[163] = 8'b01111000;
        font437[164] = 8'b11111000;
        font437[165] = 8'b01110000;
        font437[166] = 8'b00000000;
        font437[167] = 8'b00000000;
        font437[168] = 8'b00000000;
        font437[169] = 8'b01111111;
        font437[170] = 8'b01100011;
        font437[171] = 8'b01111111;
        font437[172] = 8'b01100011;
        font437[173] = 8'b01100011;
        font437[174] = 8'b01100011;
        font437[175] = 8'b01100111;
        font437[176] = 8'b11100111;
        font437[177] = 8'b11100110;
        font437[178] = 8'b11000000;
        font437[179] = 8'b00000000;
        font437[180] = 8'b00000000;
        font437[181] = 8'b00000000;
        font437[182] = 8'b00011000;
        font437[183] = 8'b11011011;
        font437[184] = 8'b01111110;
        font437[185] = 8'b11100111;
        font437[186] = 8'b11100111;
        font437[187] = 8'b01111110;
        font437[188] = 8'b11011011;
        font437[189] = 8'b00011000;
        font437[190] = 8'b00000000;
        font437[191] = 8'b00000000;
        font437[192] = 8'b00000000;
        font437[193] = 8'b10000000;
        font437[194] = 8'b11000000;
        font437[195] = 8'b11100000;
        font437[196] = 8'b11111000;
        font437[197] = 8'b11111110;
        font437[198] = 8'b11111000;
        font437[199] = 8'b11100000;
        font437[200] = 8'b11000000;
        font437[201] = 8'b10000000;
        font437[202] = 8'b00000000;
        font437[203] = 8'b00000000;
        font437[204] = 8'b00000000;
        font437[205] = 8'b00000010;
        font437[206] = 8'b00000110;
        font437[207] = 8'b00001110;
        font437[208] = 8'b00111110;
        font437[209] = 8'b11111110;
        font437[210] = 8'b00111110;
        font437[211] = 8'b00001110;
        font437[212] = 8'b00000110;
        font437[213] = 8'b00000010;
        font437[214] = 8'b00000000;
        font437[215] = 8'b00000000;
        font437[216] = 8'b00000000;
        font437[217] = 8'b00011000;
        font437[218] = 8'b00111100;
        font437[219] = 8'b01111110;
        font437[220] = 8'b00011000;
        font437[221] = 8'b00011000;
        font437[222] = 8'b00011000;
        font437[223] = 8'b01111110;
        font437[224] = 8'b00111100;
        font437[225] = 8'b00011000;
        font437[226] = 8'b00000000;
        font437[227] = 8'b00000000;
        font437[228] = 8'b00000000;
        font437[229] = 8'b01100110;
        font437[230] = 8'b01100110;
        font437[231] = 8'b01100110;
        font437[232] = 8'b01100110;
        font437[233] = 8'b01100110;
        font437[234] = 8'b00000000;
        font437[235] = 8'b00000000;
        font437[236] = 8'b01100110;
        font437[237] = 8'b01100110;
        font437[238] = 8'b00000000;
        font437[239] = 8'b00000000;
        font437[240] = 8'b00000000;
        font437[241] = 8'b01111111;
        font437[242] = 8'b11011011;
        font437[243] = 8'b11011011;
        font437[244] = 8'b11011011;
        font437[245] = 8'b01111011;
        font437[246] = 8'b00011011;
        font437[247] = 8'b00011011;
        font437[248] = 8'b00011011;
        font437[249] = 8'b00011011;
        font437[250] = 8'b00000000;
        font437[251] = 8'b00000000;
        font437[252] = 8'b00000000;
        font437[253] = 8'b01111110;
        font437[254] = 8'b01100011;
        font437[255] = 8'b00110000;
        font437[256] = 8'b00111100;
        font437[257] = 8'b01100110;
        font437[258] = 8'b01100110;
        font437[259] = 8'b00111100;
        font437[260] = 8'b00001100;
        font437[261] = 8'b11000110;
        font437[262] = 8'b01111110;
        font437[263] = 8'b00000000;
        font437[264] = 8'b00000000;
        font437[265] = 8'b00000000;
        font437[266] = 8'b00000000;
        font437[267] = 8'b00000000;
        font437[268] = 8'b00000000;
        font437[269] = 8'b00000000;
        font437[270] = 8'b00000000;
        font437[271] = 8'b11111110;
        font437[272] = 8'b11111110;
        font437[273] = 8'b11111110;
        font437[274] = 8'b00000000;
        font437[275] = 8'b00000000;
        font437[276] = 8'b00000000;
        font437[277] = 8'b00011000;
        font437[278] = 8'b00111100;
        font437[279] = 8'b01111110;
        font437[280] = 8'b00011000;
        font437[281] = 8'b00011000;
        font437[282] = 8'b00011000;
        font437[283] = 8'b01111110;
        font437[284] = 8'b00111100;
        font437[285] = 8'b00011000;
        font437[286] = 8'b01111110;
        font437[287] = 8'b00000000;
        font437[288] = 8'b00000000;
        font437[289] = 8'b00011000;
        font437[290] = 8'b00111100;
        font437[291] = 8'b01111110;
        font437[292] = 8'b00011000;
        font437[293] = 8'b00011000;
        font437[294] = 8'b00011000;
        font437[295] = 8'b00011000;
        font437[296] = 8'b00011000;
        font437[297] = 8'b00011000;
        font437[298] = 8'b00000000;
        font437[299] = 8'b00000000;
        font437[300] = 8'b00000000;
        font437[301] = 8'b00011000;
        font437[302] = 8'b00011000;
        font437[303] = 8'b00011000;
        font437[304] = 8'b00011000;
        font437[305] = 8'b00011000;
        font437[306] = 8'b00011000;
        font437[307] = 8'b01111110;
        font437[308] = 8'b00111100;
        font437[309] = 8'b00011000;
        font437[310] = 8'b00000000;
        font437[311] = 8'b00000000;
        font437[312] = 8'b00000000;
        font437[313] = 8'b00000000;
        font437[314] = 8'b00000000;
        font437[315] = 8'b00011000;
        font437[316] = 8'b00001100;
        font437[317] = 8'b11111110;
        font437[318] = 8'b00001100;
        font437[319] = 8'b00011000;
        font437[320] = 8'b00000000;
        font437[321] = 8'b00000000;
        font437[322] = 8'b00000000;
        font437[323] = 8'b00000000;
        font437[324] = 8'b00000000;
        font437[325] = 8'b00000000;
        font437[326] = 8'b00000000;
        font437[327] = 8'b00110000;
        font437[328] = 8'b01100000;
        font437[329] = 8'b11111110;
        font437[330] = 8'b01100000;
        font437[331] = 8'b00110000;
        font437[332] = 8'b00000000;
        font437[333] = 8'b00000000;
        font437[334] = 8'b00000000;
        font437[335] = 8'b00000000;
        font437[336] = 8'b00000000;
        font437[337] = 8'b00000000;
        font437[338] = 8'b00000000;
        font437[339] = 8'b00000000;
        font437[340] = 8'b11000000;
        font437[341] = 8'b11000000;
        font437[342] = 8'b11000000;
        font437[343] = 8'b11111110;
        font437[344] = 8'b00000000;
        font437[345] = 8'b00000000;
        font437[346] = 8'b00000000;
        font437[347] = 8'b00000000;
        font437[348] = 8'b00000000;
        font437[349] = 8'b00000000;
        font437[350] = 8'b00000000;
        font437[351] = 8'b00100100;
        font437[352] = 8'b01100110;
        font437[353] = 8'b11111111;
        font437[354] = 8'b01100110;
        font437[355] = 8'b00100100;
        font437[356] = 8'b00000000;
        font437[357] = 8'b00000000;
        font437[358] = 8'b00000000;
        font437[359] = 8'b00000000;
        font437[360] = 8'b00000000;
        font437[361] = 8'b00000000;
        font437[362] = 8'b00010000;
        font437[363] = 8'b00010000;
        font437[364] = 8'b00111000;
        font437[365] = 8'b00111000;
        font437[366] = 8'b01111100;
        font437[367] = 8'b01111100;
        font437[368] = 8'b11111110;
        font437[369] = 8'b11111110;
        font437[370] = 8'b00000000;
        font437[371] = 8'b00000000;
        font437[372] = 8'b00000000;
        font437[373] = 8'b00000000;
        font437[374] = 8'b11111110;
        font437[375] = 8'b11111110;
        font437[376] = 8'b01111100;
        font437[377] = 8'b01111100;
        font437[378] = 8'b00111000;
        font437[379] = 8'b00111000;
        font437[380] = 8'b00010000;
        font437[381] = 8'b00010000;
        font437[382] = 8'b00000000;
        font437[383] = 8'b00000000;
        font437[384] = 8'b00000000;
        font437[385] = 8'b00000000;
        font437[386] = 8'b00000000;
        font437[387] = 8'b00000000;
        font437[388] = 8'b00000000;
        font437[389] = 8'b00000000;
        font437[390] = 8'b00000000;
        font437[391] = 8'b00000000;
        font437[392] = 8'b00000000;
        font437[393] = 8'b00000000;
        font437[394] = 8'b00000000;
        font437[395] = 8'b00000000;
        font437[396] = 8'b00000000;
        font437[397] = 8'b00110000;
        font437[398] = 8'b01111000;
        font437[399] = 8'b01111000;
        font437[400] = 8'b01111000;
        font437[401] = 8'b00110000;
        font437[402] = 8'b00110000;
        font437[403] = 8'b00000000;
        font437[404] = 8'b00110000;
        font437[405] = 8'b00110000;
        font437[406] = 8'b00000000;
        font437[407] = 8'b00000000;
        font437[408] = 8'b00000000;
        font437[409] = 8'b01100110;
        font437[410] = 8'b01100110;
        font437[411] = 8'b01100110;
        font437[412] = 8'b00100100;
        font437[413] = 8'b00000000;
        font437[414] = 8'b00000000;
        font437[415] = 8'b00000000;
        font437[416] = 8'b00000000;
        font437[417] = 8'b00000000;
        font437[418] = 8'b00000000;
        font437[419] = 8'b00000000;
        font437[420] = 8'b00000000;
        font437[421] = 8'b01101100;
        font437[422] = 8'b01101100;
        font437[423] = 8'b11111110;
        font437[424] = 8'b01101100;
        font437[425] = 8'b01101100;
        font437[426] = 8'b01101100;
        font437[427] = 8'b11111110;
        font437[428] = 8'b01101100;
        font437[429] = 8'b01101100;
        font437[430] = 8'b00000000;
        font437[431] = 8'b00000000;
        font437[432] = 8'b00110000;
        font437[433] = 8'b00110000;
        font437[434] = 8'b01111100;
        font437[435] = 8'b11000000;
        font437[436] = 8'b11000000;
        font437[437] = 8'b01111000;
        font437[438] = 8'b00001100;
        font437[439] = 8'b00001100;
        font437[440] = 8'b11111000;
        font437[441] = 8'b00110000;
        font437[442] = 8'b00110000;
        font437[443] = 8'b00000000;
        font437[444] = 8'b00000000;
        font437[445] = 8'b00000000;
        font437[446] = 8'b00000000;
        font437[447] = 8'b11000100;
        font437[448] = 8'b11001100;
        font437[449] = 8'b00011000;
        font437[450] = 8'b00110000;
        font437[451] = 8'b01100000;
        font437[452] = 8'b11001100;
        font437[453] = 8'b10001100;
        font437[454] = 8'b00000000;
        font437[455] = 8'b00000000;
        font437[456] = 8'b00000000;
        font437[457] = 8'b01110000;
        font437[458] = 8'b11011000;
        font437[459] = 8'b11011000;
        font437[460] = 8'b01110000;
        font437[461] = 8'b11111010;
        font437[462] = 8'b11011110;
        font437[463] = 8'b11001100;
        font437[464] = 8'b11011100;
        font437[465] = 8'b01110110;
        font437[466] = 8'b00000000;
        font437[467] = 8'b00000000;
        font437[468] = 8'b00000000;
        font437[469] = 8'b00110000;
        font437[470] = 8'b00110000;
        font437[471] = 8'b00110000;
        font437[472] = 8'b01100000;
        font437[473] = 8'b00000000;
        font437[474] = 8'b00000000;
        font437[475] = 8'b00000000;
        font437[476] = 8'b00000000;
        font437[477] = 8'b00000000;
        font437[478] = 8'b00000000;
        font437[479] = 8'b00000000;
        font437[480] = 8'b00000000;
        font437[481] = 8'b00001100;
        font437[482] = 8'b00011000;
        font437[483] = 8'b00110000;
        font437[484] = 8'b01100000;
        font437[485] = 8'b01100000;
        font437[486] = 8'b01100000;
        font437[487] = 8'b00110000;
        font437[488] = 8'b00011000;
        font437[489] = 8'b00001100;
        font437[490] = 8'b00000000;
        font437[491] = 8'b00000000;
        font437[492] = 8'b00000000;
        font437[493] = 8'b01100000;
        font437[494] = 8'b00110000;
        font437[495] = 8'b00011000;
        font437[496] = 8'b00001100;
        font437[497] = 8'b00001100;
        font437[498] = 8'b00001100;
        font437[499] = 8'b00011000;
        font437[500] = 8'b00110000;
        font437[501] = 8'b01100000;
        font437[502] = 8'b00000000;
        font437[503] = 8'b00000000;
        font437[504] = 8'b00000000;
        font437[505] = 8'b00000000;
        font437[506] = 8'b00000000;
        font437[507] = 8'b01100110;
        font437[508] = 8'b00111100;
        font437[509] = 8'b11111111;
        font437[510] = 8'b00111100;
        font437[511] = 8'b01100110;
        font437[512] = 8'b00000000;
        font437[513] = 8'b00000000;
        font437[514] = 8'b00000000;
        font437[515] = 8'b00000000;
        font437[516] = 8'b00000000;
        font437[517] = 8'b00000000;
        font437[518] = 8'b00000000;
        font437[519] = 8'b00011000;
        font437[520] = 8'b00011000;
        font437[521] = 8'b01111110;
        font437[522] = 8'b00011000;
        font437[523] = 8'b00011000;
        font437[524] = 8'b00000000;
        font437[525] = 8'b00000000;
        font437[526] = 8'b00000000;
        font437[527] = 8'b00000000;
        font437[528] = 8'b00000000;
        font437[529] = 8'b00000000;
        font437[530] = 8'b00000000;
        font437[531] = 8'b00000000;
        font437[532] = 8'b00000000;
        font437[533] = 8'b00000000;
        font437[534] = 8'b00000000;
        font437[535] = 8'b00000000;
        font437[536] = 8'b00111000;
        font437[537] = 8'b00111000;
        font437[538] = 8'b01100000;
        font437[539] = 8'b00000000;
        font437[540] = 8'b00000000;
        font437[541] = 8'b00000000;
        font437[542] = 8'b00000000;
        font437[543] = 8'b00000000;
        font437[544] = 8'b00000000;
        font437[545] = 8'b11111110;
        font437[546] = 8'b00000000;
        font437[547] = 8'b00000000;
        font437[548] = 8'b00000000;
        font437[549] = 8'b00000000;
        font437[550] = 8'b00000000;
        font437[551] = 8'b00000000;
        font437[552] = 8'b00000000;
        font437[553] = 8'b00000000;
        font437[554] = 8'b00000000;
        font437[555] = 8'b00000000;
        font437[556] = 8'b00000000;
        font437[557] = 8'b00000000;
        font437[558] = 8'b00000000;
        font437[559] = 8'b00000000;
        font437[560] = 8'b00111000;
        font437[561] = 8'b00111000;
        font437[562] = 8'b00000000;
        font437[563] = 8'b00000000;
        font437[564] = 8'b00000000;
        font437[565] = 8'b00000000;
        font437[566] = 8'b00000010;
        font437[567] = 8'b00000110;
        font437[568] = 8'b00001100;
        font437[569] = 8'b00011000;
        font437[570] = 8'b00110000;
        font437[571] = 8'b01100000;
        font437[572] = 8'b11000000;
        font437[573] = 8'b10000000;
        font437[574] = 8'b00000000;
        font437[575] = 8'b00000000;
        font437[576] = 8'b00000000;
        font437[577] = 8'b01111100;
        font437[578] = 8'b11000110;
        font437[579] = 8'b11001110;
        font437[580] = 8'b11011110;
        font437[581] = 8'b11010110;
        font437[582] = 8'b11110110;
        font437[583] = 8'b11100110;
        font437[584] = 8'b11000110;
        font437[585] = 8'b01111100;
        font437[586] = 8'b00000000;
        font437[587] = 8'b00000000;
        font437[588] = 8'b00000000;
        font437[589] = 8'b00010000;
        font437[590] = 8'b00110000;
        font437[591] = 8'b11110000;
        font437[592] = 8'b00110000;
        font437[593] = 8'b00110000;
        font437[594] = 8'b00110000;
        font437[595] = 8'b00110000;
        font437[596] = 8'b00110000;
        font437[597] = 8'b11111100;
        font437[598] = 8'b00000000;
        font437[599] = 8'b00000000;
        font437[600] = 8'b00000000;
        font437[601] = 8'b01111000;
        font437[602] = 8'b11001100;
        font437[603] = 8'b11001100;
        font437[604] = 8'b00001100;
        font437[605] = 8'b00011000;
        font437[606] = 8'b00110000;
        font437[607] = 8'b01100000;
        font437[608] = 8'b11001100;
        font437[609] = 8'b11111100;
        font437[610] = 8'b00000000;
        font437[611] = 8'b00000000;
        font437[612] = 8'b00000000;
        font437[613] = 8'b01111000;
        font437[614] = 8'b11001100;
        font437[615] = 8'b00001100;
        font437[616] = 8'b00001100;
        font437[617] = 8'b00111000;
        font437[618] = 8'b00001100;
        font437[619] = 8'b00001100;
        font437[620] = 8'b11001100;
        font437[621] = 8'b01111000;
        font437[622] = 8'b00000000;
        font437[623] = 8'b00000000;
        font437[624] = 8'b00000000;
        font437[625] = 8'b00001100;
        font437[626] = 8'b00011100;
        font437[627] = 8'b00111100;
        font437[628] = 8'b01101100;
        font437[629] = 8'b11001100;
        font437[630] = 8'b11111110;
        font437[631] = 8'b00001100;
        font437[632] = 8'b00001100;
        font437[633] = 8'b00011110;
        font437[634] = 8'b00000000;
        font437[635] = 8'b00000000;
        font437[636] = 8'b00000000;
        font437[637] = 8'b11111100;
        font437[638] = 8'b11000000;
        font437[639] = 8'b11000000;
        font437[640] = 8'b11000000;
        font437[641] = 8'b11111000;
        font437[642] = 8'b00001100;
        font437[643] = 8'b00001100;
        font437[644] = 8'b11001100;
        font437[645] = 8'b01111000;
        font437[646] = 8'b00000000;
        font437[647] = 8'b00000000;
        font437[648] = 8'b00000000;
        font437[649] = 8'b00111000;
        font437[650] = 8'b01100000;
        font437[651] = 8'b11000000;
        font437[652] = 8'b11000000;
        font437[653] = 8'b11111000;
        font437[654] = 8'b11001100;
        font437[655] = 8'b11001100;
        font437[656] = 8'b11001100;
        font437[657] = 8'b01111000;
        font437[658] = 8'b00000000;
        font437[659] = 8'b00000000;
        font437[660] = 8'b00000000;
        font437[661] = 8'b11111110;
        font437[662] = 8'b11000110;
        font437[663] = 8'b11000110;
        font437[664] = 8'b00000110;
        font437[665] = 8'b00001100;
        font437[666] = 8'b00011000;
        font437[667] = 8'b00110000;
        font437[668] = 8'b00110000;
        font437[669] = 8'b00110000;
        font437[670] = 8'b00000000;
        font437[671] = 8'b00000000;
        font437[672] = 8'b00000000;
        font437[673] = 8'b01111000;
        font437[674] = 8'b11001100;
        font437[675] = 8'b11001100;
        font437[676] = 8'b11101100;
        font437[677] = 8'b01111000;
        font437[678] = 8'b11011100;
        font437[679] = 8'b11001100;
        font437[680] = 8'b11001100;
        font437[681] = 8'b01111000;
        font437[682] = 8'b00000000;
        font437[683] = 8'b00000000;
        font437[684] = 8'b00000000;
        font437[685] = 8'b01111000;
        font437[686] = 8'b11001100;
        font437[687] = 8'b11001100;
        font437[688] = 8'b11001100;
        font437[689] = 8'b01111100;
        font437[690] = 8'b00011000;
        font437[691] = 8'b00011000;
        font437[692] = 8'b00110000;
        font437[693] = 8'b01110000;
        font437[694] = 8'b00000000;
        font437[695] = 8'b00000000;
        font437[696] = 8'b00000000;
        font437[697] = 8'b00000000;
        font437[698] = 8'b00000000;
        font437[699] = 8'b00111000;
        font437[700] = 8'b00111000;
        font437[701] = 8'b00000000;
        font437[702] = 8'b00000000;
        font437[703] = 8'b00111000;
        font437[704] = 8'b00111000;
        font437[705] = 8'b00000000;
        font437[706] = 8'b00000000;
        font437[707] = 8'b00000000;
        font437[708] = 8'b00000000;
        font437[709] = 8'b00000000;
        font437[710] = 8'b00000000;
        font437[711] = 8'b00111000;
        font437[712] = 8'b00111000;
        font437[713] = 8'b00000000;
        font437[714] = 8'b00000000;
        font437[715] = 8'b00111000;
        font437[716] = 8'b00111000;
        font437[717] = 8'b00011000;
        font437[718] = 8'b00110000;
        font437[719] = 8'b00000000;
        font437[720] = 8'b00000000;
        font437[721] = 8'b00001100;
        font437[722] = 8'b00011000;
        font437[723] = 8'b00110000;
        font437[724] = 8'b01100000;
        font437[725] = 8'b11000000;
        font437[726] = 8'b01100000;
        font437[727] = 8'b00110000;
        font437[728] = 8'b00011000;
        font437[729] = 8'b00001100;
        font437[730] = 8'b00000000;
        font437[731] = 8'b00000000;
        font437[732] = 8'b00000000;
        font437[733] = 8'b00000000;
        font437[734] = 8'b00000000;
        font437[735] = 8'b00000000;
        font437[736] = 8'b01111110;
        font437[737] = 8'b00000000;
        font437[738] = 8'b01111110;
        font437[739] = 8'b00000000;
        font437[740] = 8'b00000000;
        font437[741] = 8'b00000000;
        font437[742] = 8'b00000000;
        font437[743] = 8'b00000000;
        font437[744] = 8'b00000000;
        font437[745] = 8'b01100000;
        font437[746] = 8'b00110000;
        font437[747] = 8'b00011000;
        font437[748] = 8'b00001100;
        font437[749] = 8'b00000110;
        font437[750] = 8'b00001100;
        font437[751] = 8'b00011000;
        font437[752] = 8'b00110000;
        font437[753] = 8'b01100000;
        font437[754] = 8'b00000000;
        font437[755] = 8'b00000000;
        font437[756] = 8'b00000000;
        font437[757] = 8'b01111000;
        font437[758] = 8'b11001100;
        font437[759] = 8'b00001100;
        font437[760] = 8'b00011000;
        font437[761] = 8'b00110000;
        font437[762] = 8'b00110000;
        font437[763] = 8'b00000000;
        font437[764] = 8'b00110000;
        font437[765] = 8'b00110000;
        font437[766] = 8'b00000000;
        font437[767] = 8'b00000000;
        font437[768] = 8'b00000000;
        font437[769] = 8'b01111100;
        font437[770] = 8'b11000110;
        font437[771] = 8'b11000110;
        font437[772] = 8'b11011110;
        font437[773] = 8'b11011110;
        font437[774] = 8'b11011110;
        font437[775] = 8'b11000000;
        font437[776] = 8'b11000000;
        font437[777] = 8'b01111100;
        font437[778] = 8'b00000000;
        font437[779] = 8'b00000000;
        font437[780] = 8'b00000000;
        font437[781] = 8'b00110000;
        font437[782] = 8'b01111000;
        font437[783] = 8'b11001100;
        font437[784] = 8'b11001100;
        font437[785] = 8'b11001100;
        font437[786] = 8'b11111100;
        font437[787] = 8'b11001100;
        font437[788] = 8'b11001100;
        font437[789] = 8'b11001100;
        font437[790] = 8'b00000000;
        font437[791] = 8'b00000000;
        font437[792] = 8'b00000000;
        font437[793] = 8'b11111100;
        font437[794] = 8'b01100110;
        font437[795] = 8'b01100110;
        font437[796] = 8'b01100110;
        font437[797] = 8'b01111100;
        font437[798] = 8'b01100110;
        font437[799] = 8'b01100110;
        font437[800] = 8'b01100110;
        font437[801] = 8'b11111100;
        font437[802] = 8'b00000000;
        font437[803] = 8'b00000000;
        font437[804] = 8'b00000000;
        font437[805] = 8'b00111100;
        font437[806] = 8'b01100110;
        font437[807] = 8'b11000110;
        font437[808] = 8'b11000000;
        font437[809] = 8'b11000000;
        font437[810] = 8'b11000000;
        font437[811] = 8'b11000110;
        font437[812] = 8'b01100110;
        font437[813] = 8'b00111100;
        font437[814] = 8'b00000000;
        font437[815] = 8'b00000000;
        font437[816] = 8'b00000000;
        font437[817] = 8'b11111000;
        font437[818] = 8'b01101100;
        font437[819] = 8'b01100110;
        font437[820] = 8'b01100110;
        font437[821] = 8'b01100110;
        font437[822] = 8'b01100110;
        font437[823] = 8'b01100110;
        font437[824] = 8'b01101100;
        font437[825] = 8'b11111000;
        font437[826] = 8'b00000000;
        font437[827] = 8'b00000000;
        font437[828] = 8'b00000000;
        font437[829] = 8'b11111110;
        font437[830] = 8'b01100010;
        font437[831] = 8'b01100000;
        font437[832] = 8'b01100100;
        font437[833] = 8'b01111100;
        font437[834] = 8'b01100100;
        font437[835] = 8'b01100000;
        font437[836] = 8'b01100010;
        font437[837] = 8'b11111110;
        font437[838] = 8'b00000000;
        font437[839] = 8'b00000000;
        font437[840] = 8'b00000000;
        font437[841] = 8'b11111110;
        font437[842] = 8'b01100110;
        font437[843] = 8'b01100010;
        font437[844] = 8'b01100100;
        font437[845] = 8'b01111100;
        font437[846] = 8'b01100100;
        font437[847] = 8'b01100000;
        font437[848] = 8'b01100000;
        font437[849] = 8'b11110000;
        font437[850] = 8'b00000000;
        font437[851] = 8'b00000000;
        font437[852] = 8'b00000000;
        font437[853] = 8'b00111100;
        font437[854] = 8'b01100110;
        font437[855] = 8'b11000110;
        font437[856] = 8'b11000000;
        font437[857] = 8'b11000000;
        font437[858] = 8'b11001110;
        font437[859] = 8'b11000110;
        font437[860] = 8'b01100110;
        font437[861] = 8'b00111110;
        font437[862] = 8'b00000000;
        font437[863] = 8'b00000000;
        font437[864] = 8'b00000000;
        font437[865] = 8'b11001100;
        font437[866] = 8'b11001100;
        font437[867] = 8'b11001100;
        font437[868] = 8'b11001100;
        font437[869] = 8'b11111100;
        font437[870] = 8'b11001100;
        font437[871] = 8'b11001100;
        font437[872] = 8'b11001100;
        font437[873] = 8'b11001100;
        font437[874] = 8'b00000000;
        font437[875] = 8'b00000000;
        font437[876] = 8'b00000000;
        font437[877] = 8'b01111000;
        font437[878] = 8'b00110000;
        font437[879] = 8'b00110000;
        font437[880] = 8'b00110000;
        font437[881] = 8'b00110000;
        font437[882] = 8'b00110000;
        font437[883] = 8'b00110000;
        font437[884] = 8'b00110000;
        font437[885] = 8'b01111000;
        font437[886] = 8'b00000000;
        font437[887] = 8'b00000000;
        font437[888] = 8'b00000000;
        font437[889] = 8'b00011110;
        font437[890] = 8'b00001100;
        font437[891] = 8'b00001100;
        font437[892] = 8'b00001100;
        font437[893] = 8'b00001100;
        font437[894] = 8'b11001100;
        font437[895] = 8'b11001100;
        font437[896] = 8'b11001100;
        font437[897] = 8'b01111000;
        font437[898] = 8'b00000000;
        font437[899] = 8'b00000000;
        font437[900] = 8'b00000000;
        font437[901] = 8'b11100110;
        font437[902] = 8'b01100110;
        font437[903] = 8'b01101100;
        font437[904] = 8'b01101100;
        font437[905] = 8'b01111000;
        font437[906] = 8'b01101100;
        font437[907] = 8'b01101100;
        font437[908] = 8'b01100110;
        font437[909] = 8'b11100110;
        font437[910] = 8'b00000000;
        font437[911] = 8'b00000000;
        font437[912] = 8'b00000000;
        font437[913] = 8'b11110000;
        font437[914] = 8'b01100000;
        font437[915] = 8'b01100000;
        font437[916] = 8'b01100000;
        font437[917] = 8'b01100000;
        font437[918] = 8'b01100010;
        font437[919] = 8'b01100110;
        font437[920] = 8'b01100110;
        font437[921] = 8'b11111110;
        font437[922] = 8'b00000000;
        font437[923] = 8'b00000000;
        font437[924] = 8'b00000000;
        font437[925] = 8'b11000110;
        font437[926] = 8'b11101110;
        font437[927] = 8'b11111110;
        font437[928] = 8'b11111110;
        font437[929] = 8'b11010110;
        font437[930] = 8'b11000110;
        font437[931] = 8'b11000110;
        font437[932] = 8'b11000110;
        font437[933] = 8'b11000110;
        font437[934] = 8'b00000000;
        font437[935] = 8'b00000000;
        font437[936] = 8'b00000000;
        font437[937] = 8'b11000110;
        font437[938] = 8'b11000110;
        font437[939] = 8'b11100110;
        font437[940] = 8'b11110110;
        font437[941] = 8'b11111110;
        font437[942] = 8'b11011110;
        font437[943] = 8'b11001110;
        font437[944] = 8'b11000110;
        font437[945] = 8'b11000110;
        font437[946] = 8'b00000000;
        font437[947] = 8'b00000000;
        font437[948] = 8'b00000000;
        font437[949] = 8'b00111000;
        font437[950] = 8'b01101100;
        font437[951] = 8'b11000110;
        font437[952] = 8'b11000110;
        font437[953] = 8'b11000110;
        font437[954] = 8'b11000110;
        font437[955] = 8'b11000110;
        font437[956] = 8'b01101100;
        font437[957] = 8'b00111000;
        font437[958] = 8'b00000000;
        font437[959] = 8'b00000000;
        font437[960] = 8'b00000000;
        font437[961] = 8'b11111100;
        font437[962] = 8'b01100110;
        font437[963] = 8'b01100110;
        font437[964] = 8'b01100110;
        font437[965] = 8'b01111100;
        font437[966] = 8'b01100000;
        font437[967] = 8'b01100000;
        font437[968] = 8'b01100000;
        font437[969] = 8'b11110000;
        font437[970] = 8'b00000000;
        font437[971] = 8'b00000000;
        font437[972] = 8'b00000000;
        font437[973] = 8'b00111000;
        font437[974] = 8'b01101100;
        font437[975] = 8'b11000110;
        font437[976] = 8'b11000110;
        font437[977] = 8'b11000110;
        font437[978] = 8'b11001110;
        font437[979] = 8'b11011110;
        font437[980] = 8'b01111100;
        font437[981] = 8'b00001100;
        font437[982] = 8'b00011110;
        font437[983] = 8'b00000000;
        font437[984] = 8'b00000000;
        font437[985] = 8'b11111100;
        font437[986] = 8'b01100110;
        font437[987] = 8'b01100110;
        font437[988] = 8'b01100110;
        font437[989] = 8'b01111100;
        font437[990] = 8'b01101100;
        font437[991] = 8'b01100110;
        font437[992] = 8'b01100110;
        font437[993] = 8'b11100110;
        font437[994] = 8'b00000000;
        font437[995] = 8'b00000000;
        font437[996] = 8'b00000000;
        font437[997] = 8'b01111000;
        font437[998] = 8'b11001100;
        font437[999] = 8'b11001100;
        font437[1000] = 8'b11000000;
        font437[1001] = 8'b01110000;
        font437[1002] = 8'b00011000;
        font437[1003] = 8'b11001100;
        font437[1004] = 8'b11001100;
        font437[1005] = 8'b01111000;
        font437[1006] = 8'b00000000;
        font437[1007] = 8'b00000000;
        font437[1008] = 8'b00000000;
        font437[1009] = 8'b11111100;
        font437[1010] = 8'b10110100;
        font437[1011] = 8'b00110000;
        font437[1012] = 8'b00110000;
        font437[1013] = 8'b00110000;
        font437[1014] = 8'b00110000;
        font437[1015] = 8'b00110000;
        font437[1016] = 8'b00110000;
        font437[1017] = 8'b01111000;
        font437[1018] = 8'b00000000;
        font437[1019] = 8'b00000000;
        font437[1020] = 8'b00000000;
        font437[1021] = 8'b11001100;
        font437[1022] = 8'b11001100;
        font437[1023] = 8'b11001100;
        font437[1024] = 8'b11001100;
        font437[1025] = 8'b11001100;
        font437[1026] = 8'b11001100;
        font437[1027] = 8'b11001100;
        font437[1028] = 8'b11001100;
        font437[1029] = 8'b01111000;
        font437[1030] = 8'b00000000;
        font437[1031] = 8'b00000000;
        font437[1032] = 8'b00000000;
        font437[1033] = 8'b11001100;
        font437[1034] = 8'b11001100;
        font437[1035] = 8'b11001100;
        font437[1036] = 8'b11001100;
        font437[1037] = 8'b11001100;
        font437[1038] = 8'b11001100;
        font437[1039] = 8'b11001100;
        font437[1040] = 8'b01111000;
        font437[1041] = 8'b00110000;
        font437[1042] = 8'b00000000;
        font437[1043] = 8'b00000000;
        font437[1044] = 8'b00000000;
        font437[1045] = 8'b11000110;
        font437[1046] = 8'b11000110;
        font437[1047] = 8'b11000110;
        font437[1048] = 8'b11000110;
        font437[1049] = 8'b11010110;
        font437[1050] = 8'b11010110;
        font437[1051] = 8'b01101100;
        font437[1052] = 8'b01101100;
        font437[1053] = 8'b01101100;
        font437[1054] = 8'b00000000;
        font437[1055] = 8'b00000000;
        font437[1056] = 8'b00000000;
        font437[1057] = 8'b11001100;
        font437[1058] = 8'b11001100;
        font437[1059] = 8'b11001100;
        font437[1060] = 8'b01111000;
        font437[1061] = 8'b00110000;
        font437[1062] = 8'b01111000;
        font437[1063] = 8'b11001100;
        font437[1064] = 8'b11001100;
        font437[1065] = 8'b11001100;
        font437[1066] = 8'b00000000;
        font437[1067] = 8'b00000000;
        font437[1068] = 8'b00000000;
        font437[1069] = 8'b11001100;
        font437[1070] = 8'b11001100;
        font437[1071] = 8'b11001100;
        font437[1072] = 8'b11001100;
        font437[1073] = 8'b01111000;
        font437[1074] = 8'b00110000;
        font437[1075] = 8'b00110000;
        font437[1076] = 8'b00110000;
        font437[1077] = 8'b01111000;
        font437[1078] = 8'b00000000;
        font437[1079] = 8'b00000000;
        font437[1080] = 8'b00000000;
        font437[1081] = 8'b11111110;
        font437[1082] = 8'b11001110;
        font437[1083] = 8'b10011000;
        font437[1084] = 8'b00011000;
        font437[1085] = 8'b00110000;
        font437[1086] = 8'b01100000;
        font437[1087] = 8'b01100010;
        font437[1088] = 8'b11000110;
        font437[1089] = 8'b11111110;
        font437[1090] = 8'b00000000;
        font437[1091] = 8'b00000000;
        font437[1092] = 8'b00000000;
        font437[1093] = 8'b00111100;
        font437[1094] = 8'b00110000;
        font437[1095] = 8'b00110000;
        font437[1096] = 8'b00110000;
        font437[1097] = 8'b00110000;
        font437[1098] = 8'b00110000;
        font437[1099] = 8'b00110000;
        font437[1100] = 8'b00110000;
        font437[1101] = 8'b00111100;
        font437[1102] = 8'b00000000;
        font437[1103] = 8'b00000000;
        font437[1104] = 8'b00000000;
        font437[1105] = 8'b00000000;
        font437[1106] = 8'b10000000;
        font437[1107] = 8'b11000000;
        font437[1108] = 8'b01100000;
        font437[1109] = 8'b00110000;
        font437[1110] = 8'b00011000;
        font437[1111] = 8'b00001100;
        font437[1112] = 8'b00000110;
        font437[1113] = 8'b00000010;
        font437[1114] = 8'b00000000;
        font437[1115] = 8'b00000000;
        font437[1116] = 8'b00000000;
        font437[1117] = 8'b00111100;
        font437[1118] = 8'b00001100;
        font437[1119] = 8'b00001100;
        font437[1120] = 8'b00001100;
        font437[1121] = 8'b00001100;
        font437[1122] = 8'b00001100;
        font437[1123] = 8'b00001100;
        font437[1124] = 8'b00001100;
        font437[1125] = 8'b00111100;
        font437[1126] = 8'b00000000;
        font437[1127] = 8'b00000000;
        font437[1128] = 8'b00010000;
        font437[1129] = 8'b00111000;
        font437[1130] = 8'b01101100;
        font437[1131] = 8'b11000110;
        font437[1132] = 8'b00000000;
        font437[1133] = 8'b00000000;
        font437[1134] = 8'b00000000;
        font437[1135] = 8'b00000000;
        font437[1136] = 8'b00000000;
        font437[1137] = 8'b00000000;
        font437[1138] = 8'b00000000;
        font437[1139] = 8'b00000000;
        font437[1140] = 8'b00000000;
        font437[1141] = 8'b00000000;
        font437[1142] = 8'b00000000;
        font437[1143] = 8'b00000000;
        font437[1144] = 8'b00000000;
        font437[1145] = 8'b00000000;
        font437[1146] = 8'b00000000;
        font437[1147] = 8'b00000000;
        font437[1148] = 8'b00000000;
        font437[1149] = 8'b00000000;
        font437[1150] = 8'b11111111;
        font437[1151] = 8'b00000000;
        font437[1152] = 8'b00110000;
        font437[1153] = 8'b00110000;
        font437[1154] = 8'b00011000;
        font437[1155] = 8'b00000000;
        font437[1156] = 8'b00000000;
        font437[1157] = 8'b00000000;
        font437[1158] = 8'b00000000;
        font437[1159] = 8'b00000000;
        font437[1160] = 8'b00000000;
        font437[1161] = 8'b00000000;
        font437[1162] = 8'b00000000;
        font437[1163] = 8'b00000000;
        font437[1164] = 8'b00000000;
        font437[1165] = 8'b00000000;
        font437[1166] = 8'b00000000;
        font437[1167] = 8'b00000000;
        font437[1168] = 8'b01111000;
        font437[1169] = 8'b00001100;
        font437[1170] = 8'b01111100;
        font437[1171] = 8'b11001100;
        font437[1172] = 8'b11001100;
        font437[1173] = 8'b01110110;
        font437[1174] = 8'b00000000;
        font437[1175] = 8'b00000000;
        font437[1176] = 8'b00000000;
        font437[1177] = 8'b11100000;
        font437[1178] = 8'b01100000;
        font437[1179] = 8'b01100000;
        font437[1180] = 8'b01111100;
        font437[1181] = 8'b01100110;
        font437[1182] = 8'b01100110;
        font437[1183] = 8'b01100110;
        font437[1184] = 8'b01100110;
        font437[1185] = 8'b11011100;
        font437[1186] = 8'b00000000;
        font437[1187] = 8'b00000000;
        font437[1188] = 8'b00000000;
        font437[1189] = 8'b00000000;
        font437[1190] = 8'b00000000;
        font437[1191] = 8'b00000000;
        font437[1192] = 8'b01111000;
        font437[1193] = 8'b11001100;
        font437[1194] = 8'b11000000;
        font437[1195] = 8'b11000000;
        font437[1196] = 8'b11001100;
        font437[1197] = 8'b01111000;
        font437[1198] = 8'b00000000;
        font437[1199] = 8'b00000000;
        font437[1200] = 8'b00000000;
        font437[1201] = 8'b00011100;
        font437[1202] = 8'b00001100;
        font437[1203] = 8'b00001100;
        font437[1204] = 8'b01111100;
        font437[1205] = 8'b11001100;
        font437[1206] = 8'b11001100;
        font437[1207] = 8'b11001100;
        font437[1208] = 8'b11001100;
        font437[1209] = 8'b01110110;
        font437[1210] = 8'b00000000;
        font437[1211] = 8'b00000000;
        font437[1212] = 8'b00000000;
        font437[1213] = 8'b00000000;
        font437[1214] = 8'b00000000;
        font437[1215] = 8'b00000000;
        font437[1216] = 8'b01111000;
        font437[1217] = 8'b11001100;
        font437[1218] = 8'b11111100;
        font437[1219] = 8'b11000000;
        font437[1220] = 8'b11001100;
        font437[1221] = 8'b01111000;
        font437[1222] = 8'b00000000;
        font437[1223] = 8'b00000000;
        font437[1224] = 8'b00000000;
        font437[1225] = 8'b00111000;
        font437[1226] = 8'b01101100;
        font437[1227] = 8'b01100000;
        font437[1228] = 8'b01100000;
        font437[1229] = 8'b11111000;
        font437[1230] = 8'b01100000;
        font437[1231] = 8'b01100000;
        font437[1232] = 8'b01100000;
        font437[1233] = 8'b11110000;
        font437[1234] = 8'b00000000;
        font437[1235] = 8'b00000000;
        font437[1236] = 8'b00000000;
        font437[1237] = 8'b00000000;
        font437[1238] = 8'b00000000;
        font437[1239] = 8'b00000000;
        font437[1240] = 8'b01110110;
        font437[1241] = 8'b11001100;
        font437[1242] = 8'b11001100;
        font437[1243] = 8'b11001100;
        font437[1244] = 8'b01111100;
        font437[1245] = 8'b00001100;
        font437[1246] = 8'b11001100;
        font437[1247] = 8'b01111000;
        font437[1248] = 8'b00000000;
        font437[1249] = 8'b11100000;
        font437[1250] = 8'b01100000;
        font437[1251] = 8'b01100000;
        font437[1252] = 8'b01101100;
        font437[1253] = 8'b01110110;
        font437[1254] = 8'b01100110;
        font437[1255] = 8'b01100110;
        font437[1256] = 8'b01100110;
        font437[1257] = 8'b11100110;
        font437[1258] = 8'b00000000;
        font437[1259] = 8'b00000000;
        font437[1260] = 8'b00000000;
        font437[1261] = 8'b00011000;
        font437[1262] = 8'b00011000;
        font437[1263] = 8'b00000000;
        font437[1264] = 8'b01111000;
        font437[1265] = 8'b00011000;
        font437[1266] = 8'b00011000;
        font437[1267] = 8'b00011000;
        font437[1268] = 8'b00011000;
        font437[1269] = 8'b01111110;
        font437[1270] = 8'b00000000;
        font437[1271] = 8'b00000000;
        font437[1272] = 8'b00000000;
        font437[1273] = 8'b00001100;
        font437[1274] = 8'b00001100;
        font437[1275] = 8'b00000000;
        font437[1276] = 8'b00111100;
        font437[1277] = 8'b00001100;
        font437[1278] = 8'b00001100;
        font437[1279] = 8'b00001100;
        font437[1280] = 8'b00001100;
        font437[1281] = 8'b11001100;
        font437[1282] = 8'b11001100;
        font437[1283] = 8'b01111000;
        font437[1284] = 8'b00000000;
        font437[1285] = 8'b11100000;
        font437[1286] = 8'b01100000;
        font437[1287] = 8'b01100000;
        font437[1288] = 8'b01100110;
        font437[1289] = 8'b01101100;
        font437[1290] = 8'b01111000;
        font437[1291] = 8'b01101100;
        font437[1292] = 8'b01100110;
        font437[1293] = 8'b11100110;
        font437[1294] = 8'b00000000;
        font437[1295] = 8'b00000000;
        font437[1296] = 8'b00000000;
        font437[1297] = 8'b01111000;
        font437[1298] = 8'b00011000;
        font437[1299] = 8'b00011000;
        font437[1300] = 8'b00011000;
        font437[1301] = 8'b00011000;
        font437[1302] = 8'b00011000;
        font437[1303] = 8'b00011000;
        font437[1304] = 8'b00011000;
        font437[1305] = 8'b01111110;
        font437[1306] = 8'b00000000;
        font437[1307] = 8'b00000000;
        font437[1308] = 8'b00000000;
        font437[1309] = 8'b00000000;
        font437[1310] = 8'b00000000;
        font437[1311] = 8'b00000000;
        font437[1312] = 8'b11111100;
        font437[1313] = 8'b11010110;
        font437[1314] = 8'b11010110;
        font437[1315] = 8'b11010110;
        font437[1316] = 8'b11010110;
        font437[1317] = 8'b11000110;
        font437[1318] = 8'b00000000;
        font437[1319] = 8'b00000000;
        font437[1320] = 8'b00000000;
        font437[1321] = 8'b00000000;
        font437[1322] = 8'b00000000;
        font437[1323] = 8'b00000000;
        font437[1324] = 8'b11111000;
        font437[1325] = 8'b11001100;
        font437[1326] = 8'b11001100;
        font437[1327] = 8'b11001100;
        font437[1328] = 8'b11001100;
        font437[1329] = 8'b11001100;
        font437[1330] = 8'b00000000;
        font437[1331] = 8'b00000000;
        font437[1332] = 8'b00000000;
        font437[1333] = 8'b00000000;
        font437[1334] = 8'b00000000;
        font437[1335] = 8'b00000000;
        font437[1336] = 8'b01111000;
        font437[1337] = 8'b11001100;
        font437[1338] = 8'b11001100;
        font437[1339] = 8'b11001100;
        font437[1340] = 8'b11001100;
        font437[1341] = 8'b01111000;
        font437[1342] = 8'b00000000;
        font437[1343] = 8'b00000000;
        font437[1344] = 8'b00000000;
        font437[1345] = 8'b00000000;
        font437[1346] = 8'b00000000;
        font437[1347] = 8'b00000000;
        font437[1348] = 8'b11011100;
        font437[1349] = 8'b01100110;
        font437[1350] = 8'b01100110;
        font437[1351] = 8'b01100110;
        font437[1352] = 8'b01100110;
        font437[1353] = 8'b01111100;
        font437[1354] = 8'b01100000;
        font437[1355] = 8'b11110000;
        font437[1356] = 8'b00000000;
        font437[1357] = 8'b00000000;
        font437[1358] = 8'b00000000;
        font437[1359] = 8'b00000000;
        font437[1360] = 8'b01110110;
        font437[1361] = 8'b11001100;
        font437[1362] = 8'b11001100;
        font437[1363] = 8'b11001100;
        font437[1364] = 8'b11001100;
        font437[1365] = 8'b01111100;
        font437[1366] = 8'b00001100;
        font437[1367] = 8'b00011110;
        font437[1368] = 8'b00000000;
        font437[1369] = 8'b00000000;
        font437[1370] = 8'b00000000;
        font437[1371] = 8'b00000000;
        font437[1372] = 8'b11101100;
        font437[1373] = 8'b01101110;
        font437[1374] = 8'b01110110;
        font437[1375] = 8'b01100000;
        font437[1376] = 8'b01100000;
        font437[1377] = 8'b11110000;
        font437[1378] = 8'b00000000;
        font437[1379] = 8'b00000000;
        font437[1380] = 8'b00000000;
        font437[1381] = 8'b00000000;
        font437[1382] = 8'b00000000;
        font437[1383] = 8'b00000000;
        font437[1384] = 8'b01111000;
        font437[1385] = 8'b11001100;
        font437[1386] = 8'b01100000;
        font437[1387] = 8'b00011000;
        font437[1388] = 8'b11001100;
        font437[1389] = 8'b01111000;
        font437[1390] = 8'b00000000;
        font437[1391] = 8'b00000000;
        font437[1392] = 8'b00000000;
        font437[1393] = 8'b00000000;
        font437[1394] = 8'b00100000;
        font437[1395] = 8'b01100000;
        font437[1396] = 8'b11111100;
        font437[1397] = 8'b01100000;
        font437[1398] = 8'b01100000;
        font437[1399] = 8'b01100000;
        font437[1400] = 8'b01101100;
        font437[1401] = 8'b00111000;
        font437[1402] = 8'b00000000;
        font437[1403] = 8'b00000000;
        font437[1404] = 8'b00000000;
        font437[1405] = 8'b00000000;
        font437[1406] = 8'b00000000;
        font437[1407] = 8'b00000000;
        font437[1408] = 8'b11001100;
        font437[1409] = 8'b11001100;
        font437[1410] = 8'b11001100;
        font437[1411] = 8'b11001100;
        font437[1412] = 8'b11001100;
        font437[1413] = 8'b01110110;
        font437[1414] = 8'b00000000;
        font437[1415] = 8'b00000000;
        font437[1416] = 8'b00000000;
        font437[1417] = 8'b00000000;
        font437[1418] = 8'b00000000;
        font437[1419] = 8'b00000000;
        font437[1420] = 8'b11001100;
        font437[1421] = 8'b11001100;
        font437[1422] = 8'b11001100;
        font437[1423] = 8'b11001100;
        font437[1424] = 8'b01111000;
        font437[1425] = 8'b00110000;
        font437[1426] = 8'b00000000;
        font437[1427] = 8'b00000000;
        font437[1428] = 8'b00000000;
        font437[1429] = 8'b00000000;
        font437[1430] = 8'b00000000;
        font437[1431] = 8'b00000000;
        font437[1432] = 8'b11000110;
        font437[1433] = 8'b11000110;
        font437[1434] = 8'b11010110;
        font437[1435] = 8'b11010110;
        font437[1436] = 8'b01101100;
        font437[1437] = 8'b01101100;
        font437[1438] = 8'b00000000;
        font437[1439] = 8'b00000000;
        font437[1440] = 8'b00000000;
        font437[1441] = 8'b00000000;
        font437[1442] = 8'b00000000;
        font437[1443] = 8'b00000000;
        font437[1444] = 8'b11000110;
        font437[1445] = 8'b01101100;
        font437[1446] = 8'b00111000;
        font437[1447] = 8'b00111000;
        font437[1448] = 8'b01101100;
        font437[1449] = 8'b11000110;
        font437[1450] = 8'b00000000;
        font437[1451] = 8'b00000000;
        font437[1452] = 8'b00000000;
        font437[1453] = 8'b00000000;
        font437[1454] = 8'b00000000;
        font437[1455] = 8'b00000000;
        font437[1456] = 8'b01100110;
        font437[1457] = 8'b01100110;
        font437[1458] = 8'b01100110;
        font437[1459] = 8'b01100110;
        font437[1460] = 8'b00111100;
        font437[1461] = 8'b00001100;
        font437[1462] = 8'b00011000;
        font437[1463] = 8'b11110000;
        font437[1464] = 8'b00000000;
        font437[1465] = 8'b00000000;
        font437[1466] = 8'b00000000;
        font437[1467] = 8'b00000000;
        font437[1468] = 8'b11111100;
        font437[1469] = 8'b10001100;
        font437[1470] = 8'b00011000;
        font437[1471] = 8'b01100000;
        font437[1472] = 8'b11000100;
        font437[1473] = 8'b11111100;
        font437[1474] = 8'b00000000;
        font437[1475] = 8'b00000000;
        font437[1476] = 8'b00000000;
        font437[1477] = 8'b00011100;
        font437[1478] = 8'b00110000;
        font437[1479] = 8'b00110000;
        font437[1480] = 8'b01100000;
        font437[1481] = 8'b11000000;
        font437[1482] = 8'b01100000;
        font437[1483] = 8'b00110000;
        font437[1484] = 8'b00110000;
        font437[1485] = 8'b00011100;
        font437[1486] = 8'b00000000;
        font437[1487] = 8'b00000000;
        font437[1488] = 8'b00000000;
        font437[1489] = 8'b00011000;
        font437[1490] = 8'b00011000;
        font437[1491] = 8'b00011000;
        font437[1492] = 8'b00011000;
        font437[1493] = 8'b00000000;
        font437[1494] = 8'b00011000;
        font437[1495] = 8'b00011000;
        font437[1496] = 8'b00011000;
        font437[1497] = 8'b00011000;
        font437[1498] = 8'b00000000;
        font437[1499] = 8'b00000000;
        font437[1500] = 8'b00000000;
        font437[1501] = 8'b11100000;
        font437[1502] = 8'b00110000;
        font437[1503] = 8'b00110000;
        font437[1504] = 8'b00011000;
        font437[1505] = 8'b00001100;
        font437[1506] = 8'b00011000;
        font437[1507] = 8'b00110000;
        font437[1508] = 8'b00110000;
        font437[1509] = 8'b11100000;
        font437[1510] = 8'b00000000;
        font437[1511] = 8'b00000000;
        font437[1512] = 8'b00000000;
        font437[1513] = 8'b01110011;
        font437[1514] = 8'b11011010;
        font437[1515] = 8'b11001110;
        font437[1516] = 8'b00000000;
        font437[1517] = 8'b00000000;
        font437[1518] = 8'b00000000;
        font437[1519] = 8'b00000000;
        font437[1520] = 8'b00000000;
        font437[1521] = 8'b00000000;
        font437[1522] = 8'b00000000;
        font437[1523] = 8'b00000000;
        font437[1524] = 8'b00000000;
        font437[1525] = 8'b00000000;
        font437[1526] = 8'b00000000;
        font437[1527] = 8'b00010000;
        font437[1528] = 8'b00111000;
        font437[1529] = 8'b01101100;
        font437[1530] = 8'b11000110;
        font437[1531] = 8'b11000110;
        font437[1532] = 8'b11111110;
        font437[1533] = 8'b00000000;
        font437[1534] = 8'b00000000;
        font437[1535] = 8'b00000000;
        font437[1536] = 8'b00000000;
        font437[1537] = 8'b01111000;
        font437[1538] = 8'b11001100;
        font437[1539] = 8'b11001100;
        font437[1540] = 8'b11000000;
        font437[1541] = 8'b11000000;
        font437[1542] = 8'b11000000;
        font437[1543] = 8'b11001100;
        font437[1544] = 8'b11001100;
        font437[1545] = 8'b01111000;
        font437[1546] = 8'b00110000;
        font437[1547] = 8'b11110000;
        font437[1548] = 8'b00000000;
        font437[1549] = 8'b11001100;
        font437[1550] = 8'b11001100;
        font437[1551] = 8'b00000000;
        font437[1552] = 8'b11001100;
        font437[1553] = 8'b11001100;
        font437[1554] = 8'b11001100;
        font437[1555] = 8'b11001100;
        font437[1556] = 8'b11001100;
        font437[1557] = 8'b01110110;
        font437[1558] = 8'b00000000;
        font437[1559] = 8'b00000000;
        font437[1560] = 8'b00001100;
        font437[1561] = 8'b00011000;
        font437[1562] = 8'b00110000;
        font437[1563] = 8'b00000000;
        font437[1564] = 8'b01111000;
        font437[1565] = 8'b11001100;
        font437[1566] = 8'b11111100;
        font437[1567] = 8'b11000000;
        font437[1568] = 8'b11001100;
        font437[1569] = 8'b01111000;
        font437[1570] = 8'b00000000;
        font437[1571] = 8'b00000000;
        font437[1572] = 8'b00110000;
        font437[1573] = 8'b01111000;
        font437[1574] = 8'b11001100;
        font437[1575] = 8'b00000000;
        font437[1576] = 8'b01111000;
        font437[1577] = 8'b00001100;
        font437[1578] = 8'b01111100;
        font437[1579] = 8'b11001100;
        font437[1580] = 8'b11001100;
        font437[1581] = 8'b01110110;
        font437[1582] = 8'b00000000;
        font437[1583] = 8'b00000000;
        font437[1584] = 8'b00000000;
        font437[1585] = 8'b11001100;
        font437[1586] = 8'b11001100;
        font437[1587] = 8'b00000000;
        font437[1588] = 8'b01111000;
        font437[1589] = 8'b00001100;
        font437[1590] = 8'b01111100;
        font437[1591] = 8'b11001100;
        font437[1592] = 8'b11001100;
        font437[1593] = 8'b01110110;
        font437[1594] = 8'b00000000;
        font437[1595] = 8'b00000000;
        font437[1596] = 8'b11000000;
        font437[1597] = 8'b01100000;
        font437[1598] = 8'b00110000;
        font437[1599] = 8'b00000000;
        font437[1600] = 8'b01111000;
        font437[1601] = 8'b00001100;
        font437[1602] = 8'b01111100;
        font437[1603] = 8'b11001100;
        font437[1604] = 8'b11001100;
        font437[1605] = 8'b01110110;
        font437[1606] = 8'b00000000;
        font437[1607] = 8'b00000000;
        font437[1608] = 8'b00111000;
        font437[1609] = 8'b01101100;
        font437[1610] = 8'b01101100;
        font437[1611] = 8'b00111000;
        font437[1612] = 8'b11111000;
        font437[1613] = 8'b00001100;
        font437[1614] = 8'b01111100;
        font437[1615] = 8'b11001100;
        font437[1616] = 8'b11001100;
        font437[1617] = 8'b01110110;
        font437[1618] = 8'b00000000;
        font437[1619] = 8'b00000000;
        font437[1620] = 8'b00000000;
        font437[1621] = 8'b00000000;
        font437[1622] = 8'b00000000;
        font437[1623] = 8'b00000000;
        font437[1624] = 8'b01111000;
        font437[1625] = 8'b11001100;
        font437[1626] = 8'b11000000;
        font437[1627] = 8'b11000000;
        font437[1628] = 8'b11001100;
        font437[1629] = 8'b01111000;
        font437[1630] = 8'b00110000;
        font437[1631] = 8'b11110000;
        font437[1632] = 8'b00110000;
        font437[1633] = 8'b01111000;
        font437[1634] = 8'b11001100;
        font437[1635] = 8'b00000000;
        font437[1636] = 8'b01111000;
        font437[1637] = 8'b11001100;
        font437[1638] = 8'b11111100;
        font437[1639] = 8'b11000000;
        font437[1640] = 8'b11000000;
        font437[1641] = 8'b01111100;
        font437[1642] = 8'b00000000;
        font437[1643] = 8'b00000000;
        font437[1644] = 8'b00000000;
        font437[1645] = 8'b11001100;
        font437[1646] = 8'b11001100;
        font437[1647] = 8'b00000000;
        font437[1648] = 8'b01111000;
        font437[1649] = 8'b11001100;
        font437[1650] = 8'b11111100;
        font437[1651] = 8'b11000000;
        font437[1652] = 8'b11000000;
        font437[1653] = 8'b01111100;
        font437[1654] = 8'b00000000;
        font437[1655] = 8'b00000000;
        font437[1656] = 8'b11000000;
        font437[1657] = 8'b01100000;
        font437[1658] = 8'b00110000;
        font437[1659] = 8'b00000000;
        font437[1660] = 8'b01111000;
        font437[1661] = 8'b11001100;
        font437[1662] = 8'b11111100;
        font437[1663] = 8'b11000000;
        font437[1664] = 8'b11000000;
        font437[1665] = 8'b01111100;
        font437[1666] = 8'b00000000;
        font437[1667] = 8'b00000000;
        font437[1668] = 8'b00000000;
        font437[1669] = 8'b01101100;
        font437[1670] = 8'b01101100;
        font437[1671] = 8'b00000000;
        font437[1672] = 8'b01111000;
        font437[1673] = 8'b00011000;
        font437[1674] = 8'b00011000;
        font437[1675] = 8'b00011000;
        font437[1676] = 8'b00011000;
        font437[1677] = 8'b01111110;
        font437[1678] = 8'b00000000;
        font437[1679] = 8'b00000000;
        font437[1680] = 8'b00010000;
        font437[1681] = 8'b00111000;
        font437[1682] = 8'b01101100;
        font437[1683] = 8'b00000000;
        font437[1684] = 8'b01111000;
        font437[1685] = 8'b00011000;
        font437[1686] = 8'b00011000;
        font437[1687] = 8'b00011000;
        font437[1688] = 8'b00011000;
        font437[1689] = 8'b01111110;
        font437[1690] = 8'b00000000;
        font437[1691] = 8'b00000000;
        font437[1692] = 8'b01100000;
        font437[1693] = 8'b00110000;
        font437[1694] = 8'b00011000;
        font437[1695] = 8'b00000000;
        font437[1696] = 8'b01111000;
        font437[1697] = 8'b00011000;
        font437[1698] = 8'b00011000;
        font437[1699] = 8'b00011000;
        font437[1700] = 8'b00011000;
        font437[1701] = 8'b01111110;
        font437[1702] = 8'b00000000;
        font437[1703] = 8'b00000000;
        font437[1704] = 8'b00000000;
        font437[1705] = 8'b11001100;
        font437[1706] = 8'b00000000;
        font437[1707] = 8'b00110000;
        font437[1708] = 8'b01111000;
        font437[1709] = 8'b11001100;
        font437[1710] = 8'b11001100;
        font437[1711] = 8'b11111100;
        font437[1712] = 8'b11001100;
        font437[1713] = 8'b11001100;
        font437[1714] = 8'b00000000;
        font437[1715] = 8'b00000000;
        font437[1716] = 8'b01111000;
        font437[1717] = 8'b11001100;
        font437[1718] = 8'b11001100;
        font437[1719] = 8'b01111000;
        font437[1720] = 8'b01111000;
        font437[1721] = 8'b11001100;
        font437[1722] = 8'b11001100;
        font437[1723] = 8'b11111100;
        font437[1724] = 8'b11001100;
        font437[1725] = 8'b11001100;
        font437[1726] = 8'b00000000;
        font437[1727] = 8'b00000000;
        font437[1728] = 8'b00001100;
        font437[1729] = 8'b00011000;
        font437[1730] = 8'b00110000;
        font437[1731] = 8'b11111100;
        font437[1732] = 8'b11000100;
        font437[1733] = 8'b11000000;
        font437[1734] = 8'b11111000;
        font437[1735] = 8'b11000000;
        font437[1736] = 8'b11000100;
        font437[1737] = 8'b11111100;
        font437[1738] = 8'b00000000;
        font437[1739] = 8'b00000000;
        font437[1740] = 8'b00000000;
        font437[1741] = 8'b00000000;
        font437[1742] = 8'b00000000;
        font437[1743] = 8'b00000000;
        font437[1744] = 8'b11111110;
        font437[1745] = 8'b00011011;
        font437[1746] = 8'b01111111;
        font437[1747] = 8'b11011000;
        font437[1748] = 8'b11011000;
        font437[1749] = 8'b11101111;
        font437[1750] = 8'b00000000;
        font437[1751] = 8'b00000000;
        font437[1752] = 8'b00000000;
        font437[1753] = 8'b00111110;
        font437[1754] = 8'b01111000;
        font437[1755] = 8'b11011000;
        font437[1756] = 8'b11011000;
        font437[1757] = 8'b11111110;
        font437[1758] = 8'b11011000;
        font437[1759] = 8'b11011000;
        font437[1760] = 8'b11011000;
        font437[1761] = 8'b11011110;
        font437[1762] = 8'b00000000;
        font437[1763] = 8'b00000000;
        font437[1764] = 8'b00110000;
        font437[1765] = 8'b01111000;
        font437[1766] = 8'b11001100;
        font437[1767] = 8'b00000000;
        font437[1768] = 8'b01111000;
        font437[1769] = 8'b11001100;
        font437[1770] = 8'b11001100;
        font437[1771] = 8'b11001100;
        font437[1772] = 8'b11001100;
        font437[1773] = 8'b01111000;
        font437[1774] = 8'b00000000;
        font437[1775] = 8'b00000000;
        font437[1776] = 8'b00000000;
        font437[1777] = 8'b11001100;
        font437[1778] = 8'b11001100;
        font437[1779] = 8'b00000000;
        font437[1780] = 8'b01111000;
        font437[1781] = 8'b11001100;
        font437[1782] = 8'b11001100;
        font437[1783] = 8'b11001100;
        font437[1784] = 8'b11001100;
        font437[1785] = 8'b01111000;
        font437[1786] = 8'b00000000;
        font437[1787] = 8'b00000000;
        font437[1788] = 8'b11000000;
        font437[1789] = 8'b01100000;
        font437[1790] = 8'b00110000;
        font437[1791] = 8'b00000000;
        font437[1792] = 8'b01111000;
        font437[1793] = 8'b11001100;
        font437[1794] = 8'b11001100;
        font437[1795] = 8'b11001100;
        font437[1796] = 8'b11001100;
        font437[1797] = 8'b01111000;
        font437[1798] = 8'b00000000;
        font437[1799] = 8'b00000000;
        font437[1800] = 8'b00110000;
        font437[1801] = 8'b01111000;
        font437[1802] = 8'b11001100;
        font437[1803] = 8'b00000000;
        font437[1804] = 8'b11001100;
        font437[1805] = 8'b11001100;
        font437[1806] = 8'b11001100;
        font437[1807] = 8'b11001100;
        font437[1808] = 8'b11001100;
        font437[1809] = 8'b01110110;
        font437[1810] = 8'b00000000;
        font437[1811] = 8'b00000000;
        font437[1812] = 8'b11000000;
        font437[1813] = 8'b01100000;
        font437[1814] = 8'b00110000;
        font437[1815] = 8'b00000000;
        font437[1816] = 8'b11001100;
        font437[1817] = 8'b11001100;
        font437[1818] = 8'b11001100;
        font437[1819] = 8'b11001100;
        font437[1820] = 8'b11001100;
        font437[1821] = 8'b01110110;
        font437[1822] = 8'b00000000;
        font437[1823] = 8'b00000000;
        font437[1824] = 8'b00000000;
        font437[1825] = 8'b01100110;
        font437[1826] = 8'b01100110;
        font437[1827] = 8'b00000000;
        font437[1828] = 8'b01100110;
        font437[1829] = 8'b01100110;
        font437[1830] = 8'b01100110;
        font437[1831] = 8'b01100110;
        font437[1832] = 8'b00111100;
        font437[1833] = 8'b00001100;
        font437[1834] = 8'b00011000;
        font437[1835] = 8'b11110000;
        font437[1836] = 8'b11001100;
        font437[1837] = 8'b00000000;
        font437[1838] = 8'b01111000;
        font437[1839] = 8'b11001100;
        font437[1840] = 8'b11001100;
        font437[1841] = 8'b11001100;
        font437[1842] = 8'b11001100;
        font437[1843] = 8'b11001100;
        font437[1844] = 8'b11001100;
        font437[1845] = 8'b01111000;
        font437[1846] = 8'b00000000;
        font437[1847] = 8'b00000000;
        font437[1848] = 8'b11001100;
        font437[1849] = 8'b00000000;
        font437[1850] = 8'b11001100;
        font437[1851] = 8'b11001100;
        font437[1852] = 8'b11001100;
        font437[1853] = 8'b11001100;
        font437[1854] = 8'b11001100;
        font437[1855] = 8'b11001100;
        font437[1856] = 8'b11001100;
        font437[1857] = 8'b01111000;
        font437[1858] = 8'b00000000;
        font437[1859] = 8'b00000000;
        font437[1860] = 8'b00000000;
        font437[1861] = 8'b00110000;
        font437[1862] = 8'b00110000;
        font437[1863] = 8'b01111000;
        font437[1864] = 8'b11001100;
        font437[1865] = 8'b11000000;
        font437[1866] = 8'b11000000;
        font437[1867] = 8'b11001100;
        font437[1868] = 8'b01111000;
        font437[1869] = 8'b00110000;
        font437[1870] = 8'b00110000;
        font437[1871] = 8'b00000000;
        font437[1872] = 8'b00111100;
        font437[1873] = 8'b01100110;
        font437[1874] = 8'b01100000;
        font437[1875] = 8'b01100000;
        font437[1876] = 8'b01100000;
        font437[1877] = 8'b11111100;
        font437[1878] = 8'b01100000;
        font437[1879] = 8'b01100000;
        font437[1880] = 8'b11000000;
        font437[1881] = 8'b11111110;
        font437[1882] = 8'b00000000;
        font437[1883] = 8'b00000000;
        font437[1884] = 8'b11001100;
        font437[1885] = 8'b11001100;
        font437[1886] = 8'b11001100;
        font437[1887] = 8'b11001100;
        font437[1888] = 8'b01111000;
        font437[1889] = 8'b11111100;
        font437[1890] = 8'b00110000;
        font437[1891] = 8'b11111100;
        font437[1892] = 8'b00110000;
        font437[1893] = 8'b00110000;
        font437[1894] = 8'b00000000;
        font437[1895] = 8'b00000000;
        font437[1896] = 8'b11110000;
        font437[1897] = 8'b10001000;
        font437[1898] = 8'b10001000;
        font437[1899] = 8'b10001000;
        font437[1900] = 8'b11110000;
        font437[1901] = 8'b10001000;
        font437[1902] = 8'b10011110;
        font437[1903] = 8'b10001100;
        font437[1904] = 8'b10001101;
        font437[1905] = 8'b10000110;
        font437[1906] = 8'b00000000;
        font437[1907] = 8'b00000000;
        font437[1908] = 8'b00001110;
        font437[1909] = 8'b00011011;
        font437[1910] = 8'b00011000;
        font437[1911] = 8'b00011000;
        font437[1912] = 8'b01111110;
        font437[1913] = 8'b00011000;
        font437[1914] = 8'b00011000;
        font437[1915] = 8'b00011000;
        font437[1916] = 8'b11011000;
        font437[1917] = 8'b01110000;
        font437[1918] = 8'b00000000;
        font437[1919] = 8'b00000000;
        font437[1920] = 8'b00001100;
        font437[1921] = 8'b00011000;
        font437[1922] = 8'b00110000;
        font437[1923] = 8'b00000000;
        font437[1924] = 8'b01111000;
        font437[1925] = 8'b00001100;
        font437[1926] = 8'b01111100;
        font437[1927] = 8'b11001100;
        font437[1928] = 8'b11001100;
        font437[1929] = 8'b01110110;
        font437[1930] = 8'b00000000;
        font437[1931] = 8'b00000000;
        font437[1932] = 8'b00001100;
        font437[1933] = 8'b00011000;
        font437[1934] = 8'b00110000;
        font437[1935] = 8'b00000000;
        font437[1936] = 8'b01111000;
        font437[1937] = 8'b00011000;
        font437[1938] = 8'b00011000;
        font437[1939] = 8'b00011000;
        font437[1940] = 8'b00011000;
        font437[1941] = 8'b01111110;
        font437[1942] = 8'b00000000;
        font437[1943] = 8'b00000000;
        font437[1944] = 8'b00001100;
        font437[1945] = 8'b00011000;
        font437[1946] = 8'b00110000;
        font437[1947] = 8'b00000000;
        font437[1948] = 8'b01111000;
        font437[1949] = 8'b11001100;
        font437[1950] = 8'b11001100;
        font437[1951] = 8'b11001100;
        font437[1952] = 8'b11001100;
        font437[1953] = 8'b01111000;
        font437[1954] = 8'b00000000;
        font437[1955] = 8'b00000000;
        font437[1956] = 8'b00001100;
        font437[1957] = 8'b00011000;
        font437[1958] = 8'b00110000;
        font437[1959] = 8'b00000000;
        font437[1960] = 8'b11001100;
        font437[1961] = 8'b11001100;
        font437[1962] = 8'b11001100;
        font437[1963] = 8'b11001100;
        font437[1964] = 8'b11001100;
        font437[1965] = 8'b01110110;
        font437[1966] = 8'b00000000;
        font437[1967] = 8'b00000000;
        font437[1968] = 8'b00000000;
        font437[1969] = 8'b01110110;
        font437[1970] = 8'b11011100;
        font437[1971] = 8'b00000000;
        font437[1972] = 8'b11111000;
        font437[1973] = 8'b11001100;
        font437[1974] = 8'b11001100;
        font437[1975] = 8'b11001100;
        font437[1976] = 8'b11001100;
        font437[1977] = 8'b11001100;
        font437[1978] = 8'b00000000;
        font437[1979] = 8'b00000000;
        font437[1980] = 8'b01110110;
        font437[1981] = 8'b11011100;
        font437[1982] = 8'b00000000;
        font437[1983] = 8'b11000110;
        font437[1984] = 8'b11100110;
        font437[1985] = 8'b11110110;
        font437[1986] = 8'b11011110;
        font437[1987] = 8'b11001110;
        font437[1988] = 8'b11000110;
        font437[1989] = 8'b11000110;
        font437[1990] = 8'b00000000;
        font437[1991] = 8'b00000000;
        font437[1992] = 8'b00000000;
        font437[1993] = 8'b01111000;
        font437[1994] = 8'b11001100;
        font437[1995] = 8'b11001100;
        font437[1996] = 8'b01111110;
        font437[1997] = 8'b00000000;
        font437[1998] = 8'b11111110;
        font437[1999] = 8'b00000000;
        font437[2000] = 8'b00000000;
        font437[2001] = 8'b00000000;
        font437[2002] = 8'b00000000;
        font437[2003] = 8'b00000000;
        font437[2004] = 8'b00000000;
        font437[2005] = 8'b01111000;
        font437[2006] = 8'b11001100;
        font437[2007] = 8'b11001100;
        font437[2008] = 8'b01111000;
        font437[2009] = 8'b00000000;
        font437[2010] = 8'b11111110;
        font437[2011] = 8'b00000000;
        font437[2012] = 8'b00000000;
        font437[2013] = 8'b00000000;
        font437[2014] = 8'b00000000;
        font437[2015] = 8'b00000000;
        font437[2016] = 8'b00000000;
        font437[2017] = 8'b00110000;
        font437[2018] = 8'b00110000;
        font437[2019] = 8'b00000000;
        font437[2020] = 8'b00110000;
        font437[2021] = 8'b01100000;
        font437[2022] = 8'b11000000;
        font437[2023] = 8'b11000000;
        font437[2024] = 8'b11001100;
        font437[2025] = 8'b01111000;
        font437[2026] = 8'b00000000;
        font437[2027] = 8'b00000000;
        font437[2028] = 8'b00000000;
        font437[2029] = 8'b00000000;
        font437[2030] = 8'b00000000;
        font437[2031] = 8'b00000000;
        font437[2032] = 8'b00000000;
        font437[2033] = 8'b11111100;
        font437[2034] = 8'b11000000;
        font437[2035] = 8'b11000000;
        font437[2036] = 8'b11000000;
        font437[2037] = 8'b00000000;
        font437[2038] = 8'b00000000;
        font437[2039] = 8'b00000000;
        font437[2040] = 8'b00000000;
        font437[2041] = 8'b00000000;
        font437[2042] = 8'b00000000;
        font437[2043] = 8'b00000000;
        font437[2044] = 8'b00000000;
        font437[2045] = 8'b11111100;
        font437[2046] = 8'b00001100;
        font437[2047] = 8'b00001100;
        font437[2048] = 8'b00001100;
        font437[2049] = 8'b00000000;
        font437[2050] = 8'b00000000;
        font437[2051] = 8'b00000000;
        font437[2052] = 8'b00000000;
        font437[2053] = 8'b01000010;
        font437[2054] = 8'b11000110;
        font437[2055] = 8'b11001100;
        font437[2056] = 8'b11011000;
        font437[2057] = 8'b00110000;
        font437[2058] = 8'b01101110;
        font437[2059] = 8'b11000011;
        font437[2060] = 8'b10000110;
        font437[2061] = 8'b00001100;
        font437[2062] = 8'b00011111;
        font437[2063] = 8'b00000000;
        font437[2064] = 8'b00000000;
        font437[2065] = 8'b01100011;
        font437[2066] = 8'b11100110;
        font437[2067] = 8'b01101100;
        font437[2068] = 8'b01111000;
        font437[2069] = 8'b00110111;
        font437[2070] = 8'b01101111;
        font437[2071] = 8'b11011011;
        font437[2072] = 8'b10110011;
        font437[2073] = 8'b00111111;
        font437[2074] = 8'b00000011;
        font437[2075] = 8'b00000000;
        font437[2076] = 8'b00000000;
        font437[2077] = 8'b00110000;
        font437[2078] = 8'b00110000;
        font437[2079] = 8'b00000000;
        font437[2080] = 8'b00110000;
        font437[2081] = 8'b00110000;
        font437[2082] = 8'b01111000;
        font437[2083] = 8'b01111000;
        font437[2084] = 8'b01111000;
        font437[2085] = 8'b00110000;
        font437[2086] = 8'b00000000;
        font437[2087] = 8'b00000000;
        font437[2088] = 8'b00000000;
        font437[2089] = 8'b00000000;
        font437[2090] = 8'b00000000;
        font437[2091] = 8'b00000000;
        font437[2092] = 8'b00110011;
        font437[2093] = 8'b01100110;
        font437[2094] = 8'b11001100;
        font437[2095] = 8'b11001100;
        font437[2096] = 8'b01100110;
        font437[2097] = 8'b00110011;
        font437[2098] = 8'b00000000;
        font437[2099] = 8'b00000000;
        font437[2100] = 8'b00000000;
        font437[2101] = 8'b00000000;
        font437[2102] = 8'b00000000;
        font437[2103] = 8'b00000000;
        font437[2104] = 8'b11001100;
        font437[2105] = 8'b01100110;
        font437[2106] = 8'b00110011;
        font437[2107] = 8'b00110011;
        font437[2108] = 8'b01100110;
        font437[2109] = 8'b11001100;
        font437[2110] = 8'b00000000;
        font437[2111] = 8'b00000000;
        font437[2112] = 8'b00100100;
        font437[2113] = 8'b10010010;
        font437[2114] = 8'b01001001;
        font437[2115] = 8'b00100100;
        font437[2116] = 8'b10010010;
        font437[2117] = 8'b01001001;
        font437[2118] = 8'b00100100;
        font437[2119] = 8'b10010010;
        font437[2120] = 8'b01001001;
        font437[2121] = 8'b00100100;
        font437[2122] = 8'b10010010;
        font437[2123] = 8'b01001001;
        font437[2124] = 8'b01010101;
        font437[2125] = 8'b10101010;
        font437[2126] = 8'b01010101;
        font437[2127] = 8'b10101010;
        font437[2128] = 8'b01010101;
        font437[2129] = 8'b10101010;
        font437[2130] = 8'b01010101;
        font437[2131] = 8'b10101010;
        font437[2132] = 8'b01010101;
        font437[2133] = 8'b10101010;
        font437[2134] = 8'b01010101;
        font437[2135] = 8'b10101010;
        font437[2136] = 8'b01101101;
        font437[2137] = 8'b11011011;
        font437[2138] = 8'b10110110;
        font437[2139] = 8'b01101101;
        font437[2140] = 8'b11011011;
        font437[2141] = 8'b10110110;
        font437[2142] = 8'b01101101;
        font437[2143] = 8'b11011011;
        font437[2144] = 8'b10110110;
        font437[2145] = 8'b01101101;
        font437[2146] = 8'b11011011;
        font437[2147] = 8'b10110110;
        font437[2148] = 8'b00011000;
        font437[2149] = 8'b00011000;
        font437[2150] = 8'b00011000;
        font437[2151] = 8'b00011000;
        font437[2152] = 8'b00011000;
        font437[2153] = 8'b00011000;
        font437[2154] = 8'b00011000;
        font437[2155] = 8'b00011000;
        font437[2156] = 8'b00011000;
        font437[2157] = 8'b00011000;
        font437[2158] = 8'b00011000;
        font437[2159] = 8'b00011000;
        font437[2160] = 8'b00011000;
        font437[2161] = 8'b00011000;
        font437[2162] = 8'b00011000;
        font437[2163] = 8'b00011000;
        font437[2164] = 8'b00011000;
        font437[2165] = 8'b11111000;
        font437[2166] = 8'b00011000;
        font437[2167] = 8'b00011000;
        font437[2168] = 8'b00011000;
        font437[2169] = 8'b00011000;
        font437[2170] = 8'b00011000;
        font437[2171] = 8'b00011000;
        font437[2172] = 8'b00011000;
        font437[2173] = 8'b00011000;
        font437[2174] = 8'b00011000;
        font437[2175] = 8'b00011000;
        font437[2176] = 8'b11111000;
        font437[2177] = 8'b00011000;
        font437[2178] = 8'b00011000;
        font437[2179] = 8'b11111000;
        font437[2180] = 8'b00011000;
        font437[2181] = 8'b00011000;
        font437[2182] = 8'b00011000;
        font437[2183] = 8'b00011000;
        font437[2184] = 8'b01100110;
        font437[2185] = 8'b01100110;
        font437[2186] = 8'b01100110;
        font437[2187] = 8'b01100110;
        font437[2188] = 8'b01100110;
        font437[2189] = 8'b11100110;
        font437[2190] = 8'b01100110;
        font437[2191] = 8'b01100110;
        font437[2192] = 8'b01100110;
        font437[2193] = 8'b01100110;
        font437[2194] = 8'b01100110;
        font437[2195] = 8'b01100110;
        font437[2196] = 8'b00000000;
        font437[2197] = 8'b00000000;
        font437[2198] = 8'b00000000;
        font437[2199] = 8'b00000000;
        font437[2200] = 8'b00000000;
        font437[2201] = 8'b11111110;
        font437[2202] = 8'b01100110;
        font437[2203] = 8'b01100110;
        font437[2204] = 8'b01100110;
        font437[2205] = 8'b01100110;
        font437[2206] = 8'b01100110;
        font437[2207] = 8'b01100110;
        font437[2208] = 8'b00000000;
        font437[2209] = 8'b00000000;
        font437[2210] = 8'b00000000;
        font437[2211] = 8'b00000000;
        font437[2212] = 8'b11111000;
        font437[2213] = 8'b00011000;
        font437[2214] = 8'b00011000;
        font437[2215] = 8'b11111000;
        font437[2216] = 8'b00011000;
        font437[2217] = 8'b00011000;
        font437[2218] = 8'b00011000;
        font437[2219] = 8'b00011000;
        font437[2220] = 8'b01100110;
        font437[2221] = 8'b01100110;
        font437[2222] = 8'b01100110;
        font437[2223] = 8'b01100110;
        font437[2224] = 8'b11100110;
        font437[2225] = 8'b00000110;
        font437[2226] = 8'b00000110;
        font437[2227] = 8'b11100110;
        font437[2228] = 8'b01100110;
        font437[2229] = 8'b01100110;
        font437[2230] = 8'b01100110;
        font437[2231] = 8'b01100110;
        font437[2232] = 8'b01100110;
        font437[2233] = 8'b01100110;
        font437[2234] = 8'b01100110;
        font437[2235] = 8'b01100110;
        font437[2236] = 8'b01100110;
        font437[2237] = 8'b01100110;
        font437[2238] = 8'b01100110;
        font437[2239] = 8'b01100110;
        font437[2240] = 8'b01100110;
        font437[2241] = 8'b01100110;
        font437[2242] = 8'b01100110;
        font437[2243] = 8'b01100110;
        font437[2244] = 8'b00000000;
        font437[2245] = 8'b00000000;
        font437[2246] = 8'b00000000;
        font437[2247] = 8'b00000000;
        font437[2248] = 8'b11111110;
        font437[2249] = 8'b00000110;
        font437[2250] = 8'b00000110;
        font437[2251] = 8'b11100110;
        font437[2252] = 8'b01100110;
        font437[2253] = 8'b01100110;
        font437[2254] = 8'b01100110;
        font437[2255] = 8'b01100110;
        font437[2256] = 8'b01100110;
        font437[2257] = 8'b01100110;
        font437[2258] = 8'b01100110;
        font437[2259] = 8'b01100110;
        font437[2260] = 8'b11100110;
        font437[2261] = 8'b00000110;
        font437[2262] = 8'b00000110;
        font437[2263] = 8'b11111110;
        font437[2264] = 8'b00000000;
        font437[2265] = 8'b00000000;
        font437[2266] = 8'b00000000;
        font437[2267] = 8'b00000000;
        font437[2268] = 8'b01100110;
        font437[2269] = 8'b01100110;
        font437[2270] = 8'b01100110;
        font437[2271] = 8'b01100110;
        font437[2272] = 8'b01100110;
        font437[2273] = 8'b11111110;
        font437[2274] = 8'b00000000;
        font437[2275] = 8'b00000000;
        font437[2276] = 8'b00000000;
        font437[2277] = 8'b00000000;
        font437[2278] = 8'b00000000;
        font437[2279] = 8'b00000000;
        font437[2280] = 8'b00011000;
        font437[2281] = 8'b00011000;
        font437[2282] = 8'b00011000;
        font437[2283] = 8'b00011000;
        font437[2284] = 8'b11111000;
        font437[2285] = 8'b00011000;
        font437[2286] = 8'b00011000;
        font437[2287] = 8'b11111000;
        font437[2288] = 8'b00000000;
        font437[2289] = 8'b00000000;
        font437[2290] = 8'b00000000;
        font437[2291] = 8'b00000000;
        font437[2292] = 8'b00000000;
        font437[2293] = 8'b00000000;
        font437[2294] = 8'b00000000;
        font437[2295] = 8'b00000000;
        font437[2296] = 8'b00000000;
        font437[2297] = 8'b11111000;
        font437[2298] = 8'b00011000;
        font437[2299] = 8'b00011000;
        font437[2300] = 8'b00011000;
        font437[2301] = 8'b00011000;
        font437[2302] = 8'b00011000;
        font437[2303] = 8'b00011000;
        font437[2304] = 8'b00011000;
        font437[2305] = 8'b00011000;
        font437[2306] = 8'b00011000;
        font437[2307] = 8'b00011000;
        font437[2308] = 8'b00011000;
        font437[2309] = 8'b00011111;
        font437[2310] = 8'b00000000;
        font437[2311] = 8'b00000000;
        font437[2312] = 8'b00000000;
        font437[2313] = 8'b00000000;
        font437[2314] = 8'b00000000;
        font437[2315] = 8'b00000000;
        font437[2316] = 8'b00011000;
        font437[2317] = 8'b00011000;
        font437[2318] = 8'b00011000;
        font437[2319] = 8'b00011000;
        font437[2320] = 8'b00011000;
        font437[2321] = 8'b11111111;
        font437[2322] = 8'b00000000;
        font437[2323] = 8'b00000000;
        font437[2324] = 8'b00000000;
        font437[2325] = 8'b00000000;
        font437[2326] = 8'b00000000;
        font437[2327] = 8'b00000000;
        font437[2328] = 8'b00000000;
        font437[2329] = 8'b00000000;
        font437[2330] = 8'b00000000;
        font437[2331] = 8'b00000000;
        font437[2332] = 8'b00000000;
        font437[2333] = 8'b11111111;
        font437[2334] = 8'b00011000;
        font437[2335] = 8'b00011000;
        font437[2336] = 8'b00011000;
        font437[2337] = 8'b00011000;
        font437[2338] = 8'b00011000;
        font437[2339] = 8'b00011000;
        font437[2340] = 8'b00011000;
        font437[2341] = 8'b00011000;
        font437[2342] = 8'b00011000;
        font437[2343] = 8'b00011000;
        font437[2344] = 8'b00011000;
        font437[2345] = 8'b00011111;
        font437[2346] = 8'b00011000;
        font437[2347] = 8'b00011000;
        font437[2348] = 8'b00011000;
        font437[2349] = 8'b00011000;
        font437[2350] = 8'b00011000;
        font437[2351] = 8'b00011000;
        font437[2352] = 8'b00000000;
        font437[2353] = 8'b00000000;
        font437[2354] = 8'b00000000;
        font437[2355] = 8'b00000000;
        font437[2356] = 8'b00000000;
        font437[2357] = 8'b11111111;
        font437[2358] = 8'b00000000;
        font437[2359] = 8'b00000000;
        font437[2360] = 8'b00000000;
        font437[2361] = 8'b00000000;
        font437[2362] = 8'b00000000;
        font437[2363] = 8'b00000000;
        font437[2364] = 8'b00011000;
        font437[2365] = 8'b00011000;
        font437[2366] = 8'b00011000;
        font437[2367] = 8'b00011000;
        font437[2368] = 8'b00011000;
        font437[2369] = 8'b11111111;
        font437[2370] = 8'b00011000;
        font437[2371] = 8'b00011000;
        font437[2372] = 8'b00011000;
        font437[2373] = 8'b00011000;
        font437[2374] = 8'b00011000;
        font437[2375] = 8'b00011000;
        font437[2376] = 8'b00011000;
        font437[2377] = 8'b00011000;
        font437[2378] = 8'b00011000;
        font437[2379] = 8'b00011000;
        font437[2380] = 8'b00011111;
        font437[2381] = 8'b00011000;
        font437[2382] = 8'b00011000;
        font437[2383] = 8'b00011111;
        font437[2384] = 8'b00011000;
        font437[2385] = 8'b00011000;
        font437[2386] = 8'b00011000;
        font437[2387] = 8'b00011000;
        font437[2388] = 8'b01100110;
        font437[2389] = 8'b01100110;
        font437[2390] = 8'b01100110;
        font437[2391] = 8'b01100110;
        font437[2392] = 8'b01100110;
        font437[2393] = 8'b01100111;
        font437[2394] = 8'b01100110;
        font437[2395] = 8'b01100110;
        font437[2396] = 8'b01100110;
        font437[2397] = 8'b01100110;
        font437[2398] = 8'b01100110;
        font437[2399] = 8'b01100110;
        font437[2400] = 8'b01100110;
        font437[2401] = 8'b01100110;
        font437[2402] = 8'b01100110;
        font437[2403] = 8'b01100110;
        font437[2404] = 8'b01100111;
        font437[2405] = 8'b01100000;
        font437[2406] = 8'b01100000;
        font437[2407] = 8'b01111111;
        font437[2408] = 8'b00000000;
        font437[2409] = 8'b00000000;
        font437[2410] = 8'b00000000;
        font437[2411] = 8'b00000000;
        font437[2412] = 8'b00000000;
        font437[2413] = 8'b00000000;
        font437[2414] = 8'b00000000;
        font437[2415] = 8'b00000000;
        font437[2416] = 8'b01111111;
        font437[2417] = 8'b01100000;
        font437[2418] = 8'b01100000;
        font437[2419] = 8'b01100111;
        font437[2420] = 8'b01100110;
        font437[2421] = 8'b01100110;
        font437[2422] = 8'b01100110;
        font437[2423] = 8'b01100110;
        font437[2424] = 8'b01100110;
        font437[2425] = 8'b01100110;
        font437[2426] = 8'b01100110;
        font437[2427] = 8'b01100110;
        font437[2428] = 8'b11100111;
        font437[2429] = 8'b00000000;
        font437[2430] = 8'b00000000;
        font437[2431] = 8'b11111111;
        font437[2432] = 8'b00000000;
        font437[2433] = 8'b00000000;
        font437[2434] = 8'b00000000;
        font437[2435] = 8'b00000000;
        font437[2436] = 8'b00000000;
        font437[2437] = 8'b00000000;
        font437[2438] = 8'b00000000;
        font437[2439] = 8'b00000000;
        font437[2440] = 8'b11111111;
        font437[2441] = 8'b00000000;
        font437[2442] = 8'b00000000;
        font437[2443] = 8'b11100111;
        font437[2444] = 8'b01100110;
        font437[2445] = 8'b01100110;
        font437[2446] = 8'b01100110;
        font437[2447] = 8'b01100110;
        font437[2448] = 8'b01100110;
        font437[2449] = 8'b01100110;
        font437[2450] = 8'b01100110;
        font437[2451] = 8'b01100110;
        font437[2452] = 8'b01100111;
        font437[2453] = 8'b01100000;
        font437[2454] = 8'b01100000;
        font437[2455] = 8'b01100111;
        font437[2456] = 8'b01100110;
        font437[2457] = 8'b01100110;
        font437[2458] = 8'b01100110;
        font437[2459] = 8'b01100110;
        font437[2460] = 8'b00000000;
        font437[2461] = 8'b00000000;
        font437[2462] = 8'b00000000;
        font437[2463] = 8'b00000000;
        font437[2464] = 8'b11111111;
        font437[2465] = 8'b00000000;
        font437[2466] = 8'b00000000;
        font437[2467] = 8'b11111111;
        font437[2468] = 8'b00000000;
        font437[2469] = 8'b00000000;
        font437[2470] = 8'b00000000;
        font437[2471] = 8'b00000000;
        font437[2472] = 8'b01100110;
        font437[2473] = 8'b01100110;
        font437[2474] = 8'b01100110;
        font437[2475] = 8'b01100110;
        font437[2476] = 8'b11100111;
        font437[2477] = 8'b00000000;
        font437[2478] = 8'b00000000;
        font437[2479] = 8'b11100111;
        font437[2480] = 8'b01100110;
        font437[2481] = 8'b01100110;
        font437[2482] = 8'b01100110;
        font437[2483] = 8'b01100110;
        font437[2484] = 8'b00011000;
        font437[2485] = 8'b00011000;
        font437[2486] = 8'b00011000;
        font437[2487] = 8'b00011000;
        font437[2488] = 8'b11111111;
        font437[2489] = 8'b00000000;
        font437[2490] = 8'b00000000;
        font437[2491] = 8'b11111111;
        font437[2492] = 8'b00000000;
        font437[2493] = 8'b00000000;
        font437[2494] = 8'b00000000;
        font437[2495] = 8'b00000000;
        font437[2496] = 8'b01100110;
        font437[2497] = 8'b01100110;
        font437[2498] = 8'b01100110;
        font437[2499] = 8'b01100110;
        font437[2500] = 8'b01100110;
        font437[2501] = 8'b11111111;
        font437[2502] = 8'b00000000;
        font437[2503] = 8'b00000000;
        font437[2504] = 8'b00000000;
        font437[2505] = 8'b00000000;
        font437[2506] = 8'b00000000;
        font437[2507] = 8'b00000000;
        font437[2508] = 8'b00000000;
        font437[2509] = 8'b00000000;
        font437[2510] = 8'b00000000;
        font437[2511] = 8'b00000000;
        font437[2512] = 8'b11111111;
        font437[2513] = 8'b00000000;
        font437[2514] = 8'b00000000;
        font437[2515] = 8'b11111111;
        font437[2516] = 8'b00011000;
        font437[2517] = 8'b00011000;
        font437[2518] = 8'b00011000;
        font437[2519] = 8'b00011000;
        font437[2520] = 8'b00000000;
        font437[2521] = 8'b00000000;
        font437[2522] = 8'b00000000;
        font437[2523] = 8'b00000000;
        font437[2524] = 8'b00000000;
        font437[2525] = 8'b11111111;
        font437[2526] = 8'b01100110;
        font437[2527] = 8'b01100110;
        font437[2528] = 8'b01100110;
        font437[2529] = 8'b01100110;
        font437[2530] = 8'b01100110;
        font437[2531] = 8'b01100110;
        font437[2532] = 8'b01100110;
        font437[2533] = 8'b01100110;
        font437[2534] = 8'b01100110;
        font437[2535] = 8'b01100110;
        font437[2536] = 8'b01100110;
        font437[2537] = 8'b01111111;
        font437[2538] = 8'b00000000;
        font437[2539] = 8'b00000000;
        font437[2540] = 8'b00000000;
        font437[2541] = 8'b00000000;
        font437[2542] = 8'b00000000;
        font437[2543] = 8'b00000000;
        font437[2544] = 8'b00011000;
        font437[2545] = 8'b00011000;
        font437[2546] = 8'b00011000;
        font437[2547] = 8'b00011000;
        font437[2548] = 8'b00011111;
        font437[2549] = 8'b00011000;
        font437[2550] = 8'b00011000;
        font437[2551] = 8'b00011111;
        font437[2552] = 8'b00000000;
        font437[2553] = 8'b00000000;
        font437[2554] = 8'b00000000;
        font437[2555] = 8'b00000000;
        font437[2556] = 8'b00000000;
        font437[2557] = 8'b00000000;
        font437[2558] = 8'b00000000;
        font437[2559] = 8'b00000000;
        font437[2560] = 8'b00011111;
        font437[2561] = 8'b00011000;
        font437[2562] = 8'b00011000;
        font437[2563] = 8'b00011111;
        font437[2564] = 8'b00011000;
        font437[2565] = 8'b00011000;
        font437[2566] = 8'b00011000;
        font437[2567] = 8'b00011000;
        font437[2568] = 8'b00000000;
        font437[2569] = 8'b00000000;
        font437[2570] = 8'b00000000;
        font437[2571] = 8'b00000000;
        font437[2572] = 8'b00000000;
        font437[2573] = 8'b01111111;
        font437[2574] = 8'b01100110;
        font437[2575] = 8'b01100110;
        font437[2576] = 8'b01100110;
        font437[2577] = 8'b01100110;
        font437[2578] = 8'b01100110;
        font437[2579] = 8'b01100110;
        font437[2580] = 8'b01100110;
        font437[2581] = 8'b01100110;
        font437[2582] = 8'b01100110;
        font437[2583] = 8'b01100110;
        font437[2584] = 8'b01100110;
        font437[2585] = 8'b11100111;
        font437[2586] = 8'b01100110;
        font437[2587] = 8'b01100110;
        font437[2588] = 8'b01100110;
        font437[2589] = 8'b01100110;
        font437[2590] = 8'b01100110;
        font437[2591] = 8'b01100110;
        font437[2592] = 8'b00011000;
        font437[2593] = 8'b00011000;
        font437[2594] = 8'b00011000;
        font437[2595] = 8'b00011000;
        font437[2596] = 8'b11111111;
        font437[2597] = 8'b00000000;
        font437[2598] = 8'b00000000;
        font437[2599] = 8'b11111111;
        font437[2600] = 8'b00011000;
        font437[2601] = 8'b00011000;
        font437[2602] = 8'b00011000;
        font437[2603] = 8'b00011000;
        font437[2604] = 8'b00011000;
        font437[2605] = 8'b00011000;
        font437[2606] = 8'b00011000;
        font437[2607] = 8'b00011000;
        font437[2608] = 8'b00011000;
        font437[2609] = 8'b11111000;
        font437[2610] = 8'b00000000;
        font437[2611] = 8'b00000000;
        font437[2612] = 8'b00000000;
        font437[2613] = 8'b00000000;
        font437[2614] = 8'b00000000;
        font437[2615] = 8'b00000000;
        font437[2616] = 8'b00000000;
        font437[2617] = 8'b00000000;
        font437[2618] = 8'b00000000;
        font437[2619] = 8'b00000000;
        font437[2620] = 8'b00000000;
        font437[2621] = 8'b00011111;
        font437[2622] = 8'b00011000;
        font437[2623] = 8'b00011000;
        font437[2624] = 8'b00011000;
        font437[2625] = 8'b00011000;
        font437[2626] = 8'b00011000;
        font437[2627] = 8'b00011000;
        font437[2628] = 8'b11111111;
        font437[2629] = 8'b11111111;
        font437[2630] = 8'b11111111;
        font437[2631] = 8'b11111111;
        font437[2632] = 8'b11111111;
        font437[2633] = 8'b11111111;
        font437[2634] = 8'b11111111;
        font437[2635] = 8'b11111111;
        font437[2636] = 8'b11111111;
        font437[2637] = 8'b11111111;
        font437[2638] = 8'b11111111;
        font437[2639] = 8'b11111111;
        font437[2640] = 8'b00000000;
        font437[2641] = 8'b00000000;
        font437[2642] = 8'b00000000;
        font437[2643] = 8'b00000000;
        font437[2644] = 8'b00000000;
        font437[2645] = 8'b00000000;
        font437[2646] = 8'b11111111;
        font437[2647] = 8'b11111111;
        font437[2648] = 8'b11111111;
        font437[2649] = 8'b11111111;
        font437[2650] = 8'b11111111;
        font437[2651] = 8'b11111111;
        font437[2652] = 8'b11110000;
        font437[2653] = 8'b11110000;
        font437[2654] = 8'b11110000;
        font437[2655] = 8'b11110000;
        font437[2656] = 8'b11110000;
        font437[2657] = 8'b11110000;
        font437[2658] = 8'b11110000;
        font437[2659] = 8'b11110000;
        font437[2660] = 8'b11110000;
        font437[2661] = 8'b11110000;
        font437[2662] = 8'b11110000;
        font437[2663] = 8'b11110000;
        font437[2664] = 8'b00001111;
        font437[2665] = 8'b00001111;
        font437[2666] = 8'b00001111;
        font437[2667] = 8'b00001111;
        font437[2668] = 8'b00001111;
        font437[2669] = 8'b00001111;
        font437[2670] = 8'b00001111;
        font437[2671] = 8'b00001111;
        font437[2672] = 8'b00001111;
        font437[2673] = 8'b00001111;
        font437[2674] = 8'b00001111;
        font437[2675] = 8'b00001111;
        font437[2676] = 8'b11111111;
        font437[2677] = 8'b11111111;
        font437[2678] = 8'b11111111;
        font437[2679] = 8'b11111111;
        font437[2680] = 8'b11111111;
        font437[2681] = 8'b11111111;
        font437[2682] = 8'b00000000;
        font437[2683] = 8'b00000000;
        font437[2684] = 8'b00000000;
        font437[2685] = 8'b00000000;
        font437[2686] = 8'b00000000;
        font437[2687] = 8'b00000000;
        font437[2688] = 8'b00000000;
        font437[2689] = 8'b00000000;
        font437[2690] = 8'b00000000;
        font437[2691] = 8'b00000000;
        font437[2692] = 8'b01110110;
        font437[2693] = 8'b11011110;
        font437[2694] = 8'b11001100;
        font437[2695] = 8'b11001100;
        font437[2696] = 8'b11011110;
        font437[2697] = 8'b01110110;
        font437[2698] = 8'b00000000;
        font437[2699] = 8'b00000000;
        font437[2700] = 8'b00000000;
        font437[2701] = 8'b01111000;
        font437[2702] = 8'b11001100;
        font437[2703] = 8'b11001100;
        font437[2704] = 8'b11011000;
        font437[2705] = 8'b11001100;
        font437[2706] = 8'b11001100;
        font437[2707] = 8'b11001100;
        font437[2708] = 8'b11111000;
        font437[2709] = 8'b11000000;
        font437[2710] = 8'b01100000;
        font437[2711] = 8'b00000000;
        font437[2712] = 8'b00000000;
        font437[2713] = 8'b11111100;
        font437[2714] = 8'b11001100;
        font437[2715] = 8'b11001100;
        font437[2716] = 8'b11000000;
        font437[2717] = 8'b11000000;
        font437[2718] = 8'b11000000;
        font437[2719] = 8'b11000000;
        font437[2720] = 8'b11000000;
        font437[2721] = 8'b11000000;
        font437[2722] = 8'b00000000;
        font437[2723] = 8'b00000000;
        font437[2724] = 8'b00000000;
        font437[2725] = 8'b11111110;
        font437[2726] = 8'b01101100;
        font437[2727] = 8'b01101100;
        font437[2728] = 8'b01101100;
        font437[2729] = 8'b01101100;
        font437[2730] = 8'b01101100;
        font437[2731] = 8'b01101100;
        font437[2732] = 8'b01101100;
        font437[2733] = 8'b01100110;
        font437[2734] = 8'b00000000;
        font437[2735] = 8'b00000000;
        font437[2736] = 8'b00000000;
        font437[2737] = 8'b11111100;
        font437[2738] = 8'b11000100;
        font437[2739] = 8'b01100100;
        font437[2740] = 8'b01100000;
        font437[2741] = 8'b00110000;
        font437[2742] = 8'b01100000;
        font437[2743] = 8'b01100100;
        font437[2744] = 8'b11000100;
        font437[2745] = 8'b11111100;
        font437[2746] = 8'b00000000;
        font437[2747] = 8'b00000000;
        font437[2748] = 8'b00000000;
        font437[2749] = 8'b00000000;
        font437[2750] = 8'b00000000;
        font437[2751] = 8'b00000000;
        font437[2752] = 8'b01111110;
        font437[2753] = 8'b11001000;
        font437[2754] = 8'b11001100;
        font437[2755] = 8'b11001100;
        font437[2756] = 8'b11001100;
        font437[2757] = 8'b01111000;
        font437[2758] = 8'b00000000;
        font437[2759] = 8'b00000000;
        font437[2760] = 8'b00000000;
        font437[2761] = 8'b00000000;
        font437[2762] = 8'b00000000;
        font437[2763] = 8'b00000000;
        font437[2764] = 8'b01100110;
        font437[2765] = 8'b01100110;
        font437[2766] = 8'b01100110;
        font437[2767] = 8'b01100110;
        font437[2768] = 8'b01100110;
        font437[2769] = 8'b01111011;
        font437[2770] = 8'b01100000;
        font437[2771] = 8'b11000000;
        font437[2772] = 8'b00000000;
        font437[2773] = 8'b00000000;
        font437[2774] = 8'b00000000;
        font437[2775] = 8'b01110110;
        font437[2776] = 8'b11011100;
        font437[2777] = 8'b00011000;
        font437[2778] = 8'b00011000;
        font437[2779] = 8'b00011000;
        font437[2780] = 8'b00011000;
        font437[2781] = 8'b00001110;
        font437[2782] = 8'b00000000;
        font437[2783] = 8'b00000000;
        font437[2784] = 8'b00000000;
        font437[2785] = 8'b11111100;
        font437[2786] = 8'b00110000;
        font437[2787] = 8'b01111000;
        font437[2788] = 8'b11001100;
        font437[2789] = 8'b11001100;
        font437[2790] = 8'b11001100;
        font437[2791] = 8'b01111000;
        font437[2792] = 8'b00110000;
        font437[2793] = 8'b11111100;
        font437[2794] = 8'b00000000;
        font437[2795] = 8'b00000000;
        font437[2796] = 8'b00000000;
        font437[2797] = 8'b01111000;
        font437[2798] = 8'b11001100;
        font437[2799] = 8'b11001100;
        font437[2800] = 8'b11001100;
        font437[2801] = 8'b11111100;
        font437[2802] = 8'b11001100;
        font437[2803] = 8'b11001100;
        font437[2804] = 8'b11001100;
        font437[2805] = 8'b01111000;
        font437[2806] = 8'b00000000;
        font437[2807] = 8'b00000000;
        font437[2808] = 8'b00000000;
        font437[2809] = 8'b01111100;
        font437[2810] = 8'b11000110;
        font437[2811] = 8'b11000110;
        font437[2812] = 8'b11000110;
        font437[2813] = 8'b11000110;
        font437[2814] = 8'b01101100;
        font437[2815] = 8'b01101100;
        font437[2816] = 8'b01101100;
        font437[2817] = 8'b11101110;
        font437[2818] = 8'b00000000;
        font437[2819] = 8'b00000000;
        font437[2820] = 8'b00000000;
        font437[2821] = 8'b00111100;
        font437[2822] = 8'b01100000;
        font437[2823] = 8'b00110000;
        font437[2824] = 8'b01111000;
        font437[2825] = 8'b11001100;
        font437[2826] = 8'b11001100;
        font437[2827] = 8'b11001100;
        font437[2828] = 8'b11001100;
        font437[2829] = 8'b01111000;
        font437[2830] = 8'b00000000;
        font437[2831] = 8'b00000000;
        font437[2832] = 8'b00000000;
        font437[2833] = 8'b00000000;
        font437[2834] = 8'b00000000;
        font437[2835] = 8'b01110110;
        font437[2836] = 8'b11011011;
        font437[2837] = 8'b11011011;
        font437[2838] = 8'b11011011;
        font437[2839] = 8'b01101110;
        font437[2840] = 8'b00000000;
        font437[2841] = 8'b00000000;
        font437[2842] = 8'b00000000;
        font437[2843] = 8'b00000000;
        font437[2844] = 8'b00000000;
        font437[2845] = 8'b00000000;
        font437[2846] = 8'b00000110;
        font437[2847] = 8'b01111100;
        font437[2848] = 8'b11011110;
        font437[2849] = 8'b11010110;
        font437[2850] = 8'b11110110;
        font437[2851] = 8'b01111100;
        font437[2852] = 8'b11000000;
        font437[2853] = 8'b00000000;
        font437[2854] = 8'b00000000;
        font437[2855] = 8'b00000000;
        font437[2856] = 8'b00000000;
        font437[2857] = 8'b00111100;
        font437[2858] = 8'b01100000;
        font437[2859] = 8'b11000000;
        font437[2860] = 8'b11000000;
        font437[2861] = 8'b11111100;
        font437[2862] = 8'b11000000;
        font437[2863] = 8'b11000000;
        font437[2864] = 8'b01100000;
        font437[2865] = 8'b00111100;
        font437[2866] = 8'b00000000;
        font437[2867] = 8'b00000000;
        font437[2868] = 8'b00000000;
        font437[2869] = 8'b00000000;
        font437[2870] = 8'b01111000;
        font437[2871] = 8'b11001100;
        font437[2872] = 8'b11001100;
        font437[2873] = 8'b11001100;
        font437[2874] = 8'b11001100;
        font437[2875] = 8'b11001100;
        font437[2876] = 8'b11001100;
        font437[2877] = 8'b11001100;
        font437[2878] = 8'b00000000;
        font437[2879] = 8'b00000000;
        font437[2880] = 8'b00000000;
        font437[2881] = 8'b00000000;
        font437[2882] = 8'b11111100;
        font437[2883] = 8'b00000000;
        font437[2884] = 8'b00000000;
        font437[2885] = 8'b11111100;
        font437[2886] = 8'b00000000;
        font437[2887] = 8'b00000000;
        font437[2888] = 8'b11111100;
        font437[2889] = 8'b00000000;
        font437[2890] = 8'b00000000;
        font437[2891] = 8'b00000000;
        font437[2892] = 8'b00000000;
        font437[2893] = 8'b00000000;
        font437[2894] = 8'b00110000;
        font437[2895] = 8'b00110000;
        font437[2896] = 8'b11111100;
        font437[2897] = 8'b00110000;
        font437[2898] = 8'b00110000;
        font437[2899] = 8'b00000000;
        font437[2900] = 8'b11111100;
        font437[2901] = 8'b00000000;
        font437[2902] = 8'b00000000;
        font437[2903] = 8'b00000000;
        font437[2904] = 8'b00000000;
        font437[2905] = 8'b01100000;
        font437[2906] = 8'b00110000;
        font437[2907] = 8'b00011000;
        font437[2908] = 8'b00011000;
        font437[2909] = 8'b00110000;
        font437[2910] = 8'b01100000;
        font437[2911] = 8'b00000000;
        font437[2912] = 8'b11111100;
        font437[2913] = 8'b00000000;
        font437[2914] = 8'b00000000;
        font437[2915] = 8'b00000000;
        font437[2916] = 8'b00000000;
        font437[2917] = 8'b00011000;
        font437[2918] = 8'b00110000;
        font437[2919] = 8'b01100000;
        font437[2920] = 8'b01100000;
        font437[2921] = 8'b00110000;
        font437[2922] = 8'b00011000;
        font437[2923] = 8'b00000000;
        font437[2924] = 8'b11111100;
        font437[2925] = 8'b00000000;
        font437[2926] = 8'b00000000;
        font437[2927] = 8'b00000000;
        font437[2928] = 8'b00000000;
        font437[2929] = 8'b00000000;
        font437[2930] = 8'b00001110;
        font437[2931] = 8'b00011011;
        font437[2932] = 8'b00011011;
        font437[2933] = 8'b00011000;
        font437[2934] = 8'b00011000;
        font437[2935] = 8'b00011000;
        font437[2936] = 8'b00011000;
        font437[2937] = 8'b00011000;
        font437[2938] = 8'b00011000;
        font437[2939] = 8'b00011000;
        font437[2940] = 8'b00011000;
        font437[2941] = 8'b00011000;
        font437[2942] = 8'b00011000;
        font437[2943] = 8'b00011000;
        font437[2944] = 8'b00011000;
        font437[2945] = 8'b00011000;
        font437[2946] = 8'b00011000;
        font437[2947] = 8'b11011000;
        font437[2948] = 8'b11011000;
        font437[2949] = 8'b01110000;
        font437[2950] = 8'b00000000;
        font437[2951] = 8'b00000000;
        font437[2952] = 8'b00000000;
        font437[2953] = 8'b00000000;
        font437[2954] = 8'b00110000;
        font437[2955] = 8'b00110000;
        font437[2956] = 8'b00000000;
        font437[2957] = 8'b11111100;
        font437[2958] = 8'b00000000;
        font437[2959] = 8'b00110000;
        font437[2960] = 8'b00110000;
        font437[2961] = 8'b00000000;
        font437[2962] = 8'b00000000;
        font437[2963] = 8'b00000000;
        font437[2964] = 8'b00000000;
        font437[2965] = 8'b00000000;
        font437[2966] = 8'b01110011;
        font437[2967] = 8'b11011011;
        font437[2968] = 8'b11001110;
        font437[2969] = 8'b00000000;
        font437[2970] = 8'b01110011;
        font437[2971] = 8'b11011011;
        font437[2972] = 8'b11001110;
        font437[2973] = 8'b00000000;
        font437[2974] = 8'b00000000;
        font437[2975] = 8'b00000000;
        font437[2976] = 8'b00000000;
        font437[2977] = 8'b00111100;
        font437[2978] = 8'b01100110;
        font437[2979] = 8'b01100110;
        font437[2980] = 8'b01100110;
        font437[2981] = 8'b00111100;
        font437[2982] = 8'b00000000;
        font437[2983] = 8'b00000000;
        font437[2984] = 8'b00000000;
        font437[2985] = 8'b00000000;
        font437[2986] = 8'b00000000;
        font437[2987] = 8'b00000000;
        font437[2988] = 8'b00000000;
        font437[2989] = 8'b00000000;
        font437[2990] = 8'b00000000;
        font437[2991] = 8'b00000000;
        font437[2992] = 8'b00011100;
        font437[2993] = 8'b00011100;
        font437[2994] = 8'b00000000;
        font437[2995] = 8'b00000000;
        font437[2996] = 8'b00000000;
        font437[2997] = 8'b00000000;
        font437[2998] = 8'b00000000;
        font437[2999] = 8'b00000000;
        font437[3000] = 8'b00000000;
        font437[3001] = 8'b00000000;
        font437[3002] = 8'b00000000;
        font437[3003] = 8'b00000000;
        font437[3004] = 8'b00000000;
        font437[3005] = 8'b00011000;
        font437[3006] = 8'b00000000;
        font437[3007] = 8'b00000000;
        font437[3008] = 8'b00000000;
        font437[3009] = 8'b00000000;
        font437[3010] = 8'b00000000;
        font437[3011] = 8'b00000000;
        font437[3012] = 8'b00000000;
        font437[3013] = 8'b00000111;
        font437[3014] = 8'b00000100;
        font437[3015] = 8'b00000100;
        font437[3016] = 8'b00000100;
        font437[3017] = 8'b01000100;
        font437[3018] = 8'b01100100;
        font437[3019] = 8'b00110100;
        font437[3020] = 8'b00011100;
        font437[3021] = 8'b00001100;
        font437[3022] = 8'b00000000;
        font437[3023] = 8'b00000000;
        font437[3024] = 8'b00000000;
        font437[3025] = 8'b11011000;
        font437[3026] = 8'b01101100;
        font437[3027] = 8'b01101100;
        font437[3028] = 8'b01101100;
        font437[3029] = 8'b01101100;
        font437[3030] = 8'b00000000;
        font437[3031] = 8'b00000000;
        font437[3032] = 8'b00000000;
        font437[3033] = 8'b00000000;
        font437[3034] = 8'b00000000;
        font437[3035] = 8'b00000000;
        font437[3036] = 8'b00000000;
        font437[3037] = 8'b01111000;
        font437[3038] = 8'b00001100;
        font437[3039] = 8'b00011000;
        font437[3040] = 8'b00110000;
        font437[3041] = 8'b01111100;
        font437[3042] = 8'b00000000;
        font437[3043] = 8'b00000000;
        font437[3044] = 8'b00000000;
        font437[3045] = 8'b00000000;
        font437[3046] = 8'b00000000;
        font437[3047] = 8'b00000000;
        font437[3048] = 8'b00000000;
        font437[3049] = 8'b00000000;
        font437[3050] = 8'b00111100;
        font437[3051] = 8'b00111100;
        font437[3052] = 8'b00111100;
        font437[3053] = 8'b00111100;
        font437[3054] = 8'b00111100;
        font437[3055] = 8'b00111100;
        font437[3056] = 8'b00111100;
        font437[3057] = 8'b00111100;
        font437[3058] = 8'b00000000;
        font437[3059] = 8'b00000000;
        font437[3060] = 8'b00000000;
        font437[3061] = 8'b00000000;
        font437[3062] = 8'b00000000;
        font437[3063] = 8'b00000000;
        font437[3064] = 8'b00000000;
        font437[3065] = 8'b00000000;
        font437[3066] = 8'b00000000;
        font437[3067] = 8'b00000000;
        font437[3068] = 8'b00000000;
        font437[3069] = 8'b00000000;
        font437[3070] = 8'b00000000;
        font437[3071] = 8'b00000000;
    end

    always @ (posedge clk) begin
        fontrow <= font437[faddr];
    end

    assign faddr = (char << 3) + (char << 2) + row;
    assign bits = fontrow;

endmodule
